spring !
vem ?
hjälp !
hoppa !
stanna !
vänta !
jag förstår .
jag ser .
jag vann !
le .
skål !
han sprang .
aldrig i livet !
är det sant ?
Jaså ?
tack .
vi försöker .
fråga Tom .
var trevlig .
kom igen .
släpp det !
hämta Tom .
ut med dig !
ut med er !
gå iväg .
han springer .
jag håller med .
jag instämmer .
det är okej .
kyss mig .
jag också .
perfekt !
visa mig .
berätta för mig .
vakna !
tvätta dig .
sluta !
lägg av !
var still .
stilla .
Ryck upp dig !
Ryck upp er !
kör vidare .
hitta Tom .
fixa det här .
laga den här .
Ducka .
stick !
Fortsätt in .
Hugg tag i Tom .
ha det så roligt .
Blidka mig .
gör mig till viljes .
skynda dig !
jag glömde .
jag förstår .
jag stannade kvar .
jag blev kvar .
jag använder det .
jag betalar .
jag är upptagen .
jag fryser .
det är okej med mig .
jag är ledig .
jag är mätt .
jag är hemma .
jag är sen .
jag är nästa .
jag är närmast i tur .
jag är varm .
det hjälper .
det är Tom .
det är roligt .
det är kul .
det är skoj .
det är skojigt .
kyss Tom .
låt det vara .
låt den vara .
lämna mig .
lämna oss .
gift dig med mig .
kan jag gå ?
var beredd .
håll dig redo .
håll dig i närheten .
stå upp .
Ställ dig upp !
Ställ er upp !
stanna kvar här .
sitt kvar .
stå kvar .
Ligg kvar .
Tom ljuger .
Tom grät .
Tom är uppe .
använd det här .
använd denna .
använd detta .
använd den här !
varna Tom .
se på mig .
titta på oss .
se på oss .
vem dog ?
vem har dött ?
vem slutade ?
vem är han ?
Skriv till mig .
Sikta . skjut !
sätt dig .
fåglar flyger .
Gud välsigne dig .
lugna ner dig .
lugna ner er .
lugna dig .
gör det nu .
gråt inte .
dö inte .
Ljug inte .
spring inte !
ursäkta mig .
glöm det .
ta tag i den där .
ta lite .
jag är kall .
jag kan springa .
jag kan åka skidor .
jag svimmade .
jag ger upp .
jag träffades .
jag blev träffad .
jag älskar det .
jag lovar .
jag såg en .
jag såg ett .
jag ska ringa .
jag ringer .
jag fixar maten .
jag överlever .
jag överlever nog .
jag är arg .
jag är vaken .
jag har tråkigt .
jag är pank .
jag är lycklig .
jag är tyst .
jag är tystlåten .
jag är redo !
jag är färdig !
jag är klar !
jag har rätt .
jag är nykter .
Förlåt .
jag är ung .
är det illa ?
det snöade .
den är sval .
den är cool .
det är mörkt .
det är rättvist .
det är okej .
det är gratis .
det är bra .
den är bra .
det är gott .
den är här .
den har kommit .
här är den .
den är enorm .
den är jättestor .
det är jättestort .
det är enormt .
det är mitt .
den är min .
det är okej .
den är vår .
det är vårt .
den är äkta .
det är äkta .
den är verklig .
det är sand .
det är dags .
tiden är inne .
det är sant .
det är sant .
håll dig nere .
håll er nere .
Behåll den här .
Behåll det här .
håll dig varm .
håll er varma .
släpp det .
låt mig gå !
släpp in mig .
vi försöker .
titta bort .
flytta på dig .
Självklart !
Självfallet !
Självklart .
allvarligt ?
Seriöst ?
Hen grät .
sitt stilla .
sitt still .
håll dig borta .
håll er borta .
stanna här .
sluta med det där .
sluta upp med det där .
ta min .
ta mitt .
tag min .
tag mitt .
tack .
det är okej .
det är lugnt .
sen då ?
sedan då ?
de simmade .
Tom grät .
Tom simmar .
Tom är fet .
Tom är arg .
Tom är ledsen .
Tom är blyg .
försök igen .
vi misslyckades .
vi glömde .
vi väntade .
vi kommer att vinna .
vi har vunnit !
hur är läget ?
vad händer ?
vem är han ?
vem vet ?
vem är hon ?
har jag fel ?
mår du bra ?
var belåten .
kom i tid .
var tålmodig .
ha tålamod .
var tålmodiga .
fåglar sjunger .
hämta mat .
hämta hjälp .
gå och hämta hjälp .
gå och hämta vin .
hämta vin .
får jag hjälpa ?
bär den här .
kolla det där .
kom ensam .
Självfallet !
absolut !
hoppa inte !
titta inte .
rör er inte !
rör dig inte !
Knuffas inte .
Sjung inte .
stanna inte .
prata inte !
tala inte .
vänta inte .
skrik inte .
Plikten kallar .
ät långsamt .
ät sakta .
Undersök det .
gå igenom den .
Granska den .
följ Tom .
följ efter Tom .
glöm Tom .
glöm honom .
Förlåt oss .
skaffa dig ett liv .
låt mig vara .
rör mig inte .
låt bli mig .
gå och tvätta dig !
Gud finns .
Gud existerar .
han är snäll .
han klarade det .
han hann .
han är schweizare .
han ljuger .
han är smart .
han är intelligent .
så tragiskt !
skynda dig tillbaka .
jag har tråkigt .
jag har rätt .
jag kan stanna .
jag får stanna .
jag kan simma .
det tvivlar jag på .
jag äter här .
jag känner mig vältränad .
jag känner mig ledsen .
jag hatar dig .
jag gillar honom .
jag gillar te .
jag tycker om te .
jag älskar henne .
jag älskar honom .
jag älskar dig .
jag älskar dej .
jag saknar dig .
jag behöver is .
jag behöver dig .
jag behöver er .
jag fick panik .
jag lovade .
jag minns .
jag kommer ihåg .
jag överlevde .
jag tror det .
jag ska kolla .
jag fixar det .
jag ska göra det .
jag gör det .
jag kommer att göra det .
jag kommer .
jag är hungrig .
jag är utvilad .
är Tom arg ?
är Tom galen ?
är den blå ?
är det blått ?
är det gratis ?
är det kärlek ?
är det dags ?
är tiden inne ?
är det sant ?
Jaså !
det händer .
det är mitt .
det är tomt .
det är blankt .
det står stilla .
det är uppfattat .
det är tydligt .
det är uppenbart .
den är tom .
det är tomt .
det är min cd @-@ skiva .
det är min cd .
jag bjuder .
det är säkrare .
det är läskigt .
den är läskig .
den glänser .
den sitter fast .
det sitter fast .
där är den .
det är där .
den är där .
gör det bara .
ta anteckningar .
håll still .
släpp honom !
låt den torka .
låt det torka .
släpp ut mig !
låt mig betala .
låt mig se .
titta på mig .
kärlek gör ont .
inga problem !
in med dig nu .
kom in nu .
skynda dig !
spring för livet !
hon log .
Sjung med .
stanna där .
ta en buss .
ta skydd !
prata med mig !
det är sorgligt .
det är trist .
de stod .
de röstade .
tiden flyger .
tiden rusar .
tiden är ute .
Tom kör .
Tom steg upp .
Tom slog mig .
Tom är ute .
Tom nickade .
Tom ringde .
Tom blinkade .
Tom betalar nog .
Tom är död .
Tom är döv .
Tom har dött .
Tom är snabb .
Tom är fri .
Tom är glad .
Tom är borta .
Tom har åkt .
Tom har gått .
Tom är här .
Tom är hemma .
Tom är skadad .
Tom har åkt .
Tom är säker .
Tom är svag .
Sväng höger .
vänta ett tag .
titta på det här .
kolla på det här .
vi är män .
vi är här .
vad är nytt ?
vem är hon ?
du lyckades !
du kan gå .
är du galen ?
är du arg ?
är ni arga ?
är du ny ?
är du ledsen ?
var kreativ .
var kreativa .
var diskret .
var diskreta .
var vänlig .
var vänliga .
var generös .
var generösa .
var nådig .
var redo .
var punktlig .
var punktliga .
var hänsynslös .
var förnuftig .
var specifik .
var tydlig .
var tolerant .
var toleranta .
var vaksam .
var vaksamma .
var på din vakt .
var på er vakt .
öl är gott .
kolla en gång till .
kom närmare .
kom in .
trösta Tom .
kontakta Tom .
ta kontakt med Tom .
vann du ?
gör det igen !
gör det igen .
gör det senare .
gör det rätt .
inga men .
Fuska inte .
gör det inte !
gör det inte .
slåss inte .
Glo inte .
gå inte .
skjut inte !
le inte .
tala inte .
prata inte .
stå inte .
Stirra inte .
oroa dig inte .
byt om .
byt kläder .
klä på dig .
klä på er .
gå och hämta hjälp .
gå med Tom .
följ med Tom .
han får komma .
han kan simma .
han ljuger .
han gillar mig .
han älskar mig .
han blev skadad .
han blev sårad .
han låtsas .
han är stark .
hur är det ?
hur mår du ?
jag gick också .
jag är längre .
jag kan köra .
jag kan inte äta .
jag äter frukt .
jag fick ett jobb .
jag skaffade mig ett jobb .
jag fastnade .
jag blev trött .
jag hatar arbete .
jag gillar båda .
jag gillar jazz .
jag gillar det här .
jag bor här .
jag älskar rock .
jag försov mig .
jag hämtade mig .
jag ordnade det .
jag säljer bilar .
jag tackar dig .
jag tackar er .
jag litar på er .
jag var arg .
jag blev avskedad .
jag hade tur .
jag var trött .
jag arbetar här .
jag jobbar här .
jag ska byta om .
jag klarar mig .
jag hämtar den .
jag hämtar det .
jag är hemma .
jag är säker .
jag är nyfiken .
jag är ursinnig .
jag är rasande .
jag är hälsosam .
jag är seriös .
jag är utsvulten .
jag är törstig .
jag är rörd .
jag vinner .
är Tom näst i tur ?
är det vitt ?
är hon trevlig ?
det hände .
det kommer kanske att göra ont .
det är måndag .
det är meningslöst .
den är låst .
det är mitt jobb .
det är normalt .
det är vanligt .
in med dig bara .
låt mig hjälpa till .
låt mig leva .
livet är roligt .
Lunchen är klar .
Lunchen är färdig .
ingen kom .
snälla kom .
snälla sluta !
hon bet honom .
hon slog honom .
hon är snäll .
stå still !
stå stilla !
stanna inomhus .
rör dig inte .
sluta försöka .
tala långsammare .
det är okej .
det där är okej .
det är bra .
Sånt är livet .
sådant är livet .
det är mitt .
det är okej .
det är sant .
tv:n är på .
de kysste varandra .
det här är dåligt .
Tom fnissade .
Tom blev biten .
Tom är tillbaka .
Tom är död .
Tom är döv .
Tom är fattig .
Tom är lång .
Tom är svag .
Tom klarade sig .
Tom lyckades .
Tom gjorde den .
Tom gjorde det .
Tom undervisar .
Tom var stor .
Tom ringer nog .
Tom kommer nog .
Tom hjälper nog till .
Tom överlever .
Tom överlever nog .
Tom tänker sluta .
Tom stannar nog .
Tom väntar nog .
Tom är alert .
Tom är på alerten .
Tom är uppmärksam .
Tom är snabb i vändningarna .
Tom är vid liv .
Tom är ensam .
Tom är allena .
Tom är för sig själv .
Tom är arg .
Tom är vaken .
Tom är uttråkad .
Tom är tokig .
Tom är galen .
Tom är full .
Tom dör .
Tom är tidig .
Tom är stollig .
Tom är hispig .
Tom är knäpp .
Tom är rolig .
Tom har tur .
Tom är lyckligt lottad .
Tom ljuger .
Tom är framfusig .
Tom är framåt .
Tom har rätt .
Tom är smart .
Tom är trött .
Tom har fel .
Tom är ung .
stäng av den .
hade jag fel ?
vi åt ägg .
vi gjorde slut .
vi behöver dig .
vi lovade .
vi överlevde .
vi är döende .
vi ska åka .
vi ska gå .
vi åker .
vi går .
vi är färdiga .
vi är klara .
vi är redo .
vad är nytt ?
vad kommer härnäst ?
vad ska ske nu ?
vad händer nu ?
vad är detta ?
var är han ?
vem flydde ?
vem går först ?
vem är först i tur ?
vem står först i tur ?
du är min .
är jag förälskad ?
är du vilse ?
är du säker ?
är du utom fara ?
är du trygg ?
är du tillräknelig ?
är du vid dina sinnens fulla bruk ?
är ni tillräkneliga ?
är ni vid era sinnens fulla bruk ?
är du säker ?
är det säkert ?
Koka ett ägg .
gå och hämta förstärkning .
kan du komma ?
kan du simma ?
kom framåt .
kom fram .
kom fort !
kom med oss .
har Tom ringt ?
röstade Tom ?
röstade du ?
ser jag OK ut ?
ser jag bra ut ?
gör det på måndag .
gör det ändå .
håller ni med ?
röker ni ?
röker du ?
Snarkar du ?
fråga inte mig .
var inte ledsen .
Skämta inte med mig !
släpp inte taget .
skrik inte .
kör fortare .
kör försiktigt .
Visitera dem .
Undersök dem .
Undersök den här .
hitta katten .
fisk , tack .
gå tillbaka , Tom .
gå dit nu .
god morgon !
Väx upp , Tom .
håll ut , Tom .
ta dig ett glas .
ta en drink .
ta en till .
han kan göra det .
han har en bil .
han har hund .
han har en hund .
han är en poet .
han äter .
han älskar henne .
han drev med mig .
han var själv .
han var ensam .
han var modig .
han var mäktig .
han var jättebra .
han kommer att komma .
han kommer att gå .
han är så söt .
hjälp mig , Tom .
hjälp oss , Tom .
vad spännande !
vad patetiskt !
hur går det på skolan ?
hur går det i skolan ?
jag är hemma .
jag är så sjuk .
jag bad om ursäkt .
jag kan försöka göra det .
jag bryr mig inte .
jag har inget emot det .
jag har en katt .
jag har ett jobb .
jag har ett barn .
jag har en penna .
jag måste gå .
jag improviserade .
jag känner till en väg .
jag vet ett sätt .
jag vet en väg .
jag gillar frukt .
jag tycker om frukt .
jag älskar att resa .
jag hittade på det .
jag stannar kanske .
jag behöver en hatt .
jag behöver ett jobb .
jag behöver en penna .
jag behöver målarfärg .
jag behövde dig .
jag behövde er .
jag ser en bok .
jag fattar .
jag förstår .
jag fattar .
jag förstår .
jag promenerar mycket .
jag går mycket .
jag var hungrig .
jag drog mig ur .
jag kommer inte att förlora .
jag flyttar inte .
jag flyttar mig inte .
jag flyttar inte på mig .
jag undrar varför .
jag klarar mig .
jag kommer att vara här .
jag är här .
jag fixar en .
jag hämtar en .
jag ska betala dig .
jag ska spara det .
jag är doktor .
jag är konstnärlig .
jag är konstnärligt lagd .
jag är konstnärlig av mig .
jag är upptagen nu .
jag drunknar .
jag flyr .
jag är färdig .
jag är hemsk .
jag har slutat med öl .
jag är så lycklig .
jag är bäst .
jag är kittlig .
det är mitt fel .
jag är jättetjock .
jag fick dig .
jag har dig .
går måndag bra ?
går det bra på måndag ?
funkar måndag ?
fungerar måndag ?
är Tom galen ?
är det sant ?
är detta kärlek ?
den var svart .
det var svart .
det var natt .
det var högljutt .
den var högljudd .
det var tyst .
den var tyst .
den var rund .
det var runt .
det är pinsamt .
den är äkta .
det är äkta .
den är autentisk .
det är autentiskt .
det haglar .
det är inget skämt .
det är konstigt .
den är konstig .
det är märkligt .
det är underligt .
den är för stor .
det är för varmt .
den fungerar .
det fungerar .
den funkar .
det funkar .
Fortsätt dansa .
Fortsätt springa .
Fortsätt le .
Fortsätt tala .
Fortsätt arbeta .
Damerna först .
låt Tom leva .
låt Tom stanna .
låt mig göra det .
Mary kom in .
det gör ont i mina öron .
behöver jag fortsätta ?
ingen vet .
ingen vet .
snälla ta det lugnt .
snälla lugna ner dig .
peka ut den .
peka ut det .
hon kan simma .
hon är lycklig .
hon är tystlåten .
hon är tyst .
hon känner mig .
hon gillade det .
hon gillade den .
hon tyckte om det .
hon tyckte om den .
hon gick ut .
tala långsammare .
stanna bilen .
det är mitt .
den är min .
vad hemskt .
det är smart .
vad konstigt .
de störtade .
de kraschlandade .
de gjorde bankrutt .
de gick i kras .
de kraschade .
de vill ha mig .
de kommer att misslyckas .
de kommer att växa .
de är blå .
de är deppiga .
de är färdiga .
de är klara .
Tom blev klar .
Tom blev färdig .
Tom lyckades fly .
Tom kom hem .
Tom tog sig hem .
Tom gick vilse .
Tom har dött .
Tom har ryggrad .
Tom har kurage .
Tom hatade det .
Tom hatade den .
Tom hatar tv .
Tom hatar mig .
Tom hörde det .
Tom hjälper oss .
Tom anställde mig .
Tom slog Mary .
Tom lever .
Tom är vaken .
Tom är hemsk .
Tom är mörkhyad .
Tom är pank .
Tom är grym .
Tom är yr .
Tom ljuger .
Tom är naiv .
Tom behöver mig .
Tom sa ja .
Tom ryckte på axlarna .
Tom var mätt .
Tom var nyfiken .
Tom är road .
Tom gråter .
Tom äter .
Tom är känd .
Tom är smutsig .
Tom är lortig .
Tom är snål .
Tom är ostadig på benen .
Tom är groggy .
Tom är skyldig .
Tom är hungrig .
Tom är mentalsjuk .
Tom är sinnessjuk .
Tom är vansinnig .
Tom skämtar .
Tom är ensam .
Tom är inte här .
Tom är inte på .
Tom är artig .
Tom är rädd .
Tom är tyst .
Tom är hög .
Tom är sträng .
Tom är stark .
vi är araber .
vi kommer överens .
vi kommer väl överens .
vi bor här .
vi måste prata .
vi måste pratas vid .
vi måste tala .
vi måste talas vid .
vi behöver hjälp .
vi klarar oss .
vi är på insidan .
vi är inne .
vi försöker .
vad är det ?
vad är detta ?
vad är det här ?
du är sen .
du är lat !
ni är lata !
du ser tjock ut .
du får stanna .
ni får stanna .
du kan stanna .
ni kan stanna .
du får simma .
du verkar ledsen .
du överlevde .
ni överlevde .
du är döende .
du ljuger !
du är konstig .
du har vuxit .
är jag säker nu ?
någonting annat ?
är du ett fan ?
är du galen ?
var respektfull .
ring snuten .
får jag fråga vem ?
får jag ta den ?
kan vi gå nu ?
kom imorgon .
gjorde jag det där ?
var det jag som gjorde det där ?
gjorde du det ?
gjorde ni det ?
känner jag Tom ?
känner jag honom ?
behöver jag en ?
drömmer katter ?
gör det genast .
gör det snabbt .
gör det fort .
gör det tyst .
fattar du ?
vet Tom ?
vet Tom om det ?
hundar kan simma .
var inte elak .
var inte oförskämd .
var inte ohövlig .
var inte ohyfsad .
gör inte det här .
gör inte detta .
ge inte upp !
var inte uppkäftig .
var inte kaxig .
rita en cirkel .
skynda på dig .
skynda på er .
Sno på dig .
Sno på er .
skynda på .
Raska på .
rör på benen .
kom hit .
hämta hjälp .
ge mig en dag .
ge mig en pistol .
ge mig ett jobb .
ge mig ett arbete .
gå och hämta en öl .
gå och hämta kaffe .
ge den till mig .
håll i den .
ta en kaka .
han drack öl .
han kände sig trött .
han har en blogg .
han kramade henne .
han är min typ !
han dödade honom .
han ljög för oss .
han ser blek ut .
han ljuger aldrig .
han verkar snäll .
han går fort .
Hen grät .
han blev blind .
han är besvärlig .
han är inget helgon .
han är inte sjuk .
han studerar .
han pluggar .
här kommer han .
han blödde näsblod .
håll fast i den .
håll i repet .
håll repet .
du då ?
hur illa är det ?
hur varm är den ?
hur varmt är det ?
hur sen är jag ?
Tom , skynda dig .
jag går alltid .
jag är i Paris .
jag åt snabbt .
jag tror på dig .
jag kan vara rättvis .
jag kan vara snäll .
jag kan vara trevlig .
jag kan köpa två .
jag kan köpa två stycken .
jag kan göra båda .
jag kan göra mer .
jag kan göra mera .
det kan jag göra .
jag kan inte dansa .
jag gjorde det som jag skulle göra .
jag gjorde ingenting .
jag gillar verkligen Tom .
jag känner mig ensam .
jag somnade .
jag föll för den .
jag var hungrig .
jag hade ingen aning .
jag var tvungen att gömma mig .
jag är förkyld .
jag har en ring .
jag har en fru .
jag lät Tom vinna .
jag ljög för Tom .
jag ljög för dig .
jag ljög för er .
jag gillar filmer .
jag tycker om filmer .
jag tycker om mitt jobb .
jag tycker om tennis .
jag gillar tåg .
jag tycker om tåg .
jag gillar vinter .
jag bor i närheten .
jag älskar arabiska .
jag älskar äpplen .
jag älskar hästar .
jag älskar min katt .
jag älskar min mamma .
jag gillar vinter .
jag gjorde upp en affär .
jag saknar Boston .
jag måste gå nu .
jag måste bege mig nu .
jag behöver en plan .
jag behöver kaffe .
jag behöver den nu .
jag måste försöka .
jag behövde det här .
jag är skyldig Tom en .
jag äger en lustjakt .
jag äger en yacht .
jag satte den tillbaka .
jag driver ett motell .
jag såg Tom dö .
jag såg ett flygplan .
jag såg honom gråta .
det ordnade jag .
det såg jag till .
jag ser mitt skepp .
jag sålde en bok .
jag berättade ett skämt .
jag använder Firefox .
jag vill ha en tårta .
jag vill ha alltsamman .
jag vill ha alltsammans .
jag vill vinna .
jag var hemma .
jag blev drogad .
jag var kär .
jag var orolig .
jag väckte dig .
jag jobbar natt .
jag går först .
jag kommer att gå först .
jag hjälper dig .
jag ska hjälpa dig .
jag kommer att hjälpa dig .
jag ska berätta för dig .
jag kommer att berätta för dig .
jag berättar för dig .
jag är man nu .
jag är vacker .
jag är också här .
jag är bara lat .
jag är motiverad .
jag är peppad .
jag är ingen expert .
jag är inte någon expert .
jag är objektiv .
jag är nöjd .
jag är belåten .
jag är för ung .
jag är väldigt upptagen .
är min tid slut ?
det kunde funka .
det är liknande .
det är likt .
den är liknande .
den är lik .
det kommer inte att fungera .
det kommer inte att funka .
det kommer inte att gå .
det är lördag .
den är övergiven .
det har hänt .
det är min häst .
det är möjligt .
det är för kallt .
den är för kall .
det är för högt .
den är väldigt stor .
Fortsätt klättra .
hör av dig !
låt honom göra det .
låt mig hämta den .
låt mig hämta det .
vi ger upp .
vi provar en .
vi testar en .
vi smakar på en .
livet är galet .
Lås dörren !
Mary är konstig .
får jag gå hem ?
mamma är på jobbet .
det värker i huvudet .
det är ingen hemma .
nu kan vi gå .
nu kan vi åka .
okej , hör på .
öppna dörren .
vårt lag förlorade .
ta det lugnt .
ta det i din egen takt .
Välj ett nummer .
säg något .
ska jag fortsätta ?
hon undviker mig .
hon böjde sig ner .
hon böjde sig ned .
hon kom sist .
hon blev arg .
hon hatade honom .
hon hatar honom .
hon hjälper honom .
hon är tvilling .
hon gråter .
hon gillar honom .
hon ser ledsen ut .
hon ser lessen ut .
hon älskar Tom .
hon älskar honom .
hon var modig .
hon gick hem .
hon åkte hem .
hon for hem .
hon är grym .
hon håller diet .
hon är min typ .
hon är min fru .
Tänk positivt .
var positiv .
se det positiva .
sluta skjuta !
sluta skjuta !
sluta oroa dig .
ta bara en .
det var svårt .
den där var enorm .
den där var vår .
det där är Saturnus .
det är en plan .
det är ju helt befängt !
det är bättre .
det är genomförbart .
det är mycket .
det är enkelt .
det är så typiskt dig .
de lämnade återbud .
de omfamnade varandra .
de älskade det .
de älskade den .
de är panka .
de är barskrapade .
de är nära .
de är unga .
det här är en penna .
det här är konstigt .
detta är konstigt .
detta är underligt .
det här är underligt .
Tom böjde sig ned .
Tom köpte den .
Tom köpte det .
Tom gick på det .
Tom gick på den .
Tom gick med på det .
Tom kom sist .
Tom gjorde bra ifrån sig .
Tom tränade .
Tom tränar .
Tom kände sig sårad .
Tom blev yr .
Tom fick sparken .
Tom blev avskedad .
Tom blev glad .
Tom har planer .
Tom har annat för sig .
Tom hatar dig .
Tom hatar er .
Tom är en sportig typ .
Tom är en idrottare .
Tom är en idrottskille .
Tom är en nörd .
Tom är en tölp .
Tom är en drummel .
Tom är en fårskalle .
Tom är en luns .
Tom är utomlands .
Tom är inte här .
Tom är frånvarande .
Tom är aktiv .
Tom är livlig .
Tom är road .
Tom är skärpt .
Tom är knubbig .
Tom är smart .
Tom är listig .
Tom är bakslug .
Tom är knäpp .
Tom är vresig .
Tom är rättfram .
Tom äter .
Tom är i min ålder .
Tom är inte rolig .
Tom är artig .
Tom är rädd .
Tom är stark .
Tom lämnade hemmet .
Tom reste hemifrån .
Tom släppte in mig .
Tom lät oss gå .
Tom tycker om dig .
Tom gillar dig .
Tom ser sjuk ut .
Tom ser gammal ut .
Tom frisknade till .
Tom tillfrisknade .
Tom springer snabbt .
Tom vill ha en .
Tom var yr .
Tom blev anställd .
Tom hade rätt .
Tom åkte tillbaka .
Tom gick tillbaka .
Tom klarar sig nog .
Tom är adopterad .
Tom är ängslig .
Tom har anlänt .
Tom håller på att kvävas .
Tom lagar mat .
Tom har rätt .
Tom är förlovad .
Tom har rymt .
Tom har svimmat .
Tom är ursinnig .
Tom hjälper till .
Tom hjälper .
Tom haltar .
Tom är gift .
Tom är inte tjock .
Tom packar .
Tom vilar .
Tom är pensionerad .
Tom är ärlig .
Tom är konstig .
Tom väntar .
Tom arbetar .
Tom är orolig .
Tom är ängslig .
Tom är bekymrad .
försök göra det .
försök att göra det .
var Tom ensam ?
vatten , tack .
vi kan få ett slut på det .
vi kan få ett slut på den .
vi kan använda det .
vi kan inte misslyckas .
vi fick punktering .
vi måste gå .
vi såg alltihop .
vi förstår .
vi vill ha fred .
vi ville ha Tom .
vi var panka .
vi hade rätt .
vi kommer att klara det .
vi kommer att överleva .
vi är oroliga .
vi är försiktiga .
vi är noggranna .
vi är noga .
vilken lättnad !
vilken relief !
vad får jag ?
vad var det som hände ?
vad ska vi göra ?
vad ska vi ta oss till ?
när var det ?
var är du ?
var är ni ?
vilken är min ?
vem hatar dig ?
Vilka är det som hatar dig ?
Vilka är det som hatar er ?
vem kör ?
vem vinner ?
varför ändra på det ?
kommer hon att komma ?
du klarar det .
du kan göra det .
det klarar du .
det klarar du av .
du ser upptagen ut .
du ser sjuk ut .
du behöver det här .
du behöver den här .
du borde gå .
du talar fort .
ni talar fort .
du talar snabbt .
ni talar snabbt .
du pratar snabbt .
ni pratar snabbt .
du är en snobb .
du är partisk .
du är inte rolig .
du är så het .
ni är så heta .
du är dum .
du är fånig .
du är orättvis .
ni är orättvisa .
är jag misstänkt ?
är vi vänner ?
sover du ?
är du partisk ?
är ni partiska ?
är du fördomsfull ?
är ni fördomsfulla ?
har ni fördomar ?
har du förutfattade meningar ?
har ni förutfattade meningar ?
gråter du ?
Grinar du ?
är du hungrig ?
är ni hungriga ?
har jag inte rätt ?
är inte du Tom ?
var snäll med Tom .
var snäll mot henne .
Fåglarna lägger ägg .
fåglar lägger ägg .
får jag vara där ?
kan jag ringa dig ?
kan jag ringa er ?
får jag också komma ?
kan jag få en ?
kan jag hjälpa dig ?
kan jag komma med dig ?
får jag träffa dem ?
får jag se dem ?
kan jag få se dem ?
kan jag få träffa dem ?
får jag också se ?
kan jag sitta ned ?
får jag tala nu ?
kan jag använda den här ?
kan vi komma in ?
kan vi göra det ?
kan vi gå hem ?
får vi behålla den ?
klarar vi det ?
kan vi flytta den ?
kan du laga den ?
kan du sitta upprätt ?
kan du sitta rak ?
städa rummet .
kom tillbaka hit .
kom och sitt bredvid mig .
kor äter gräs .
pappa är inte hemma .
det är roligt att dansa .
det är kul att dansa .
köpte Tom den ?
gick det bra ?
gjorde vi bra ifrån oss ?
hade vi det ?
klarade vi det ?
åkte ni allihopa ?
lagade du den ?
fattade du ?
provade du det ?
använde du den ?
middagen är klar !
middagen är färdig !
gör som Tom säger .
gör som du vill .
gör det nu , Tom .
gör det så här .
gör det på det här sättet .
gör det i morgon .
gör det själv .
har vi någon ?
känner vi dig ?
känner vi er ?
gillar du den ?
gillar du det ?
älskar du det ?
Älskaru mej ?
saknar du det ?
saknar du mig ?
lovar du ?
lovar ni ?
var inte arg .
var inte ohyfsad .
sluta larva dig .
Ställ dig inte upp .
rör mig inte !
titta inte på tv .
bryr du dig inte ?
ät allting .
alla ner på marken !
alla visste .
alla gick .
alla betalade .
alla flämtar .
alla är ute .
in i bilen med dig .
sätt dig i bilen .
släpp Tom .
gör dig av med Tom .
gör er av med Tom .
sov lite .
sätt igång , Tom .
ge den åt Tom .
ge den till henne .
ge den till honom .
ge det till honom .
ge mig en öl .
ge mig skjuts .
ge mig ett tecken .
ge mig en vecka .
ge mig min väska .
gå och hälsa på Tom .
gå och byt om .
gå och ta en öl .
gå och hämta Tom .
gå och prata med Tom .
Goddag .
ta dina saker .
gott nytt år !
god fortsättning !
har Tom ringt ?
har de åkt ?
har du ätit ?
han var nära att dö .
han bad mig göra det .
han kan inte simma .
han förtjänade det .
han fick jobbet .
han hade en radio .
han höll i en boll .
han är författare .
han är stilig .
han är min fiende .
han bor ensam .
han ser ung ut .
han älskar musik .
han är skyldig mig det .
det verkar som om han är trött .
han verkar trött .
det verkar som att han är trött .
han promenerade hem .
han gick hem .
han var hemma .
han var min chef .
han var törstig .
han är lite blyg .
han är lite blyg av sig .
här kommer Tom .
här är bussen .
hej , stig på .
hans huvud värkte .
han hade huvudvärk .
Bromsa .
håll den åt mig .
hur illa var det ?
hur dåligt var det ?
hur kan jag hjälpa till ?
hur kan jag hjälpa ?
hur kallt är det ?
hur gick det för dig ?
hur ska jag göra det ?
hur ser vi ut ?
hur långt borta var det ?
hur svårt är det ?
hur sent är det ?
hur var Hawaii ?
jag vet redan .
jag är i London .
jag åt en banan .
jag åt upp alla .
jag åt för mycket .
jag ringde i förväg .
jag kom för att hjälpa till .
jag kan hämta den .
jag kan höra dig .
jag kan hjälpa dig .
jag kan döda dig .
jag kan ta livet av dig .
jag kan ta Tom .
jag kan köra Tom .
jag kan bättre än sådär .
det kan jag försöka göra .
jag gjorde det igen .
jag varnade faktiskt Tom .
jag sov inte .
jag ogillar ägg .
jag menar verkligen det .
jag fattar inte .
jag dricker kaffe .
jag blev förälskad .
jag gav bort den .
jag avslöjade den .
jag återlämnade den .
jag gav den tillbaka .
jag fattar .
jag går till skolan .
jag växte upp här .
jag roade mig .
jag var tvungen att åka i väg .
jag var tvungen att åka .
jag hatar måndagar .
jag hatar Tom nu .
jag hatar den också .
jag hatar karaoke .
jag hatar min kropp .
jag hatar mitt hår .
jag hatar spindlar .
jag avskyr att stryka .
jag hatar att stryka .
jag har ett kännetecken .
jag har en bricka .
jag har ett emblem .
jag har ett märke .
jag har ett ordenstecken .
jag har feber .
jag har en flöjt .
jag har en idé .
jag har haft roligt .
jag har haft kul .
jag har inga barn .
jag har kartan .
jag måste hjälpa till .
jag måste gömma mig
jag måste vila .
jag måste stanna .
jag måste vänta .
jag hörde en duns .
jag hörde röster .
jag gjorde illa foten .
jag gjorde mig illa i foten .
jag träffade honom precis .
jag vill bara ha den .
jag skriver dagbok .
jag för dagbok .
jag gjorde Tom besviken .
jag svek Tom .
jag övergav Tom .
jag lät Tom tala .
jag tycker om att köra bil .
jag tycker om lasagne .
jag tycker om att fiska .
jag bor i norra delen av staten .
jag tappade kontrollen .
jag älskar bananer .
jag hittade på det där .
jag kan ha rätt .
jag träffade Tom här .
jag träffade honom en gång .
jag saknar min fru .
jag måste vara lugn .
jag behöver en kniv .
jag behöver en handduk .
jag behöver min jacka .
jag behöver min rock .
jag behöver min kappa .
jag behöver en nu .
jag behöver dig nu .
jag går aldrig ut .
jag såg den aldrig .
jag reser ofta .
jag betalade kontant .
jag betalade med kontanter .
jag betalar Tom bra .
jag vägrar gå .
jag sa stick .
lägg av , sa jag .
inte nu , sa jag .
håll käften , sa jag .
ta den , sa jag .
jag såg Tom falla .
jag såg henne simma .
jag såg honom en gång .
jag såg ett en gång .
jag ser boken .
jag tjänar ingen .
jag har verkligen kallt .
det hoppas jag verkligen .
jag slängde ut den .
jag tog det lugnt .
jag promenerar till jobbet .
jag vill ha fläkten .
jag vill rösta .
jag var inte i tjänst .
jag var tjänstledig .
jag sov .
det var mitt fel .
jag var för snabb .
jag kommer att få ett slut på det .
jag kommer att stoppa det .
jag tar den .
jag vann loppet .
jag arbetar för Tom .
jag skrev till Tom .
jag ska be om ursäkt .
jag hämtar Tom .
jag ska göra det nu .
jag tar hand om det .
jag kommer att sakna det .
jag betalar extra .
jag ska betala extra .
jag kommer att betala extra .
jag ska skjuta dig .
jag kommer att skjuta dig .
jag väntar här .
jag kommer att vänta här .
jag är Toms fru .
jag är musiker .
jag är pacifist .
jag är arg på dig .
jag är inte hungrig .
jag är precis här .
jag är mållös .
jag är mördaren .
jag har gjort det .
är det så illa ?
är hon hemma ?
är det där franska ?
är det här franska ?
är det här franskt ?
är det här fransk ?
den är inte billig .
den såg äkta ut .
det låter enkelt .
det gör fortfarande ont .
det var en dröm .
det var kaotiskt .
det var korrekt .
det snöade .
det är jul .
då är det avgjort .
det är ett problem .
den är ett problem .
det är svårt .
den är svår .
det är dyrt .
det är varmt i dag .
det är viktigt .
den är viktig .
det är nödvändigt .
det är meningslöst .
det är sant .
den är för liten .
det är för litet .
det går att behandla .
lämna mig ifred !
låt mig vara !
lämna mig i fred !
lämna mig ifred .
låt mig hämta Tom .
livet är orättvist .
lyssna på detta !
Lev och lär .
Lunchen är klar .
Lunchen är färdig .
Lynn springer snabbt .
många fiskar dog .
får jag kyssa dig ?
min hund bet Tom .
mitt jobb är säkert .
det värker i lederna .
jag heter Tom .
ingen skrek .
ingen berättade det för oss .
ingen blev träffad .
ingen är upprörd .
gör det nu bara .
stanna där nu .
öppna era ögon .
säg det tydligt .
vi ses på måndag .
ska vi dansa ?
ska vi beställa ?
hon kom ensam .
hon lurade honom .
hon hjälpte honom .
hon kramade honom .
hon är sjuksköterska .
hon är ute nu .
hon sparkade honom .
hon gillar vin .
hon såg ledsen ut .
hon älskar katter .
hon kommer kanske .
hon saknar honom .
hon ljuger aldrig .
hon sjunger bra .
hon simmar bra .
Hen grät .
hon är en ängel .
visa oss runt .
våren är här .
håll dig bakom mig .
håll er bakom mig .
sommaren är över .
ta tid på dig .
ta det lugnt .
ingen brådska .
Förta dig för all del inte .
det där var läskigt .
de körde fort .
det är en början .
det är min replik .
det är min fru .
det där är plast .
det är allvarligt .
det är självmord .
det är förräderi .
det var oturligt .
radion dog .
de har rätt .
de köpte det .
de köpte den .
de kan dö .
de hatade Tom .
de kramade oss .
de ser bra ut .
de bråkade .
de litar på dig .
de var mina .
de kommer inte att dö .
de kommer att attackera .
de kommer att anfalla .
de är rädda .
de har gått sönder .
det här är min väska .
detta är min bil .
det här är min bil .
de där är gratis .
de där är trevliga .
de där är fina .
biljetten , tack .
dags att stiga upp .
dags att gå upp .
Tom kan inte komma .
Tom kan inte läsa .
Tom kan inte stanna .
Tom kan inte gå .
Tom klappade ihop .
Tom tog knäcken på sig .
Tom dog ensam .
Tom dog vid 65 .
Tom kom närmare .
Tom blev dumpad .
Tom blev rädd .
Tom odlar ris .
Tom hade cancer .
Tom har utslag .
Tom har tandställning .
Tom har problem .
Tom har min bil .
Tom har talang .
Tom hatar katter .
Tom avskyr katter .
Tom hatar råttor .
Tom hörde Mary .
Tom hörde det där .
Tom anställde Mary .
Tom är ett äckel .
Tom är en haj .
Tom är en svindlare .
Tom är rolig .
Tom är orolig .
Tom är ängslig .
Tom är skamsen .
Tom är toppen .
Tom är grym .
Tom är besvärlig .
Tom är förbryllad .
Tom är säker .
Tom är oärlig .
Tom är bedräglig .
Tom är hängiven .
Tom är påklädd .
Tom är tveksam .
Tom är förlovad .
Tom är rasande .
Tom är gift .
Tom saknas .
Tom är min hjälte .
Tom är neutral .
Tom nickar .
Tom är omtyckt .
Tom är populär .
Tom väntar .
Tom arbetar .
Tom är inte död .
Tom är inte här .
Tom är inte lat .
Tom är inte trevlig .
Tom är inte fattig .
Tom är inte otrevlig .
Tom är inte smal .
Tom är inte ful .
Tom tycker om snö .
Tom gillar snö .
Tom tycker om vin .
Tom såg sjuk ut .
Tom såg gammal ut .
Tom såg ledsen ut .
Tom ser blek ut .
Tom ser illamående ut .
Tom saknar dig .
Tom behöver hjälp .
Tom tuppade av .
Tom svimmade .
Tom kolade av .
Tom dog .
Tom verkar trevlig .
Tom grät .
Tom blev rånad .
Tom kommer inte att stanna .
Tom återhämtar sig nog .
Tom kommer nog att lyckas .
Tom överlever nog .
Tom blöder .
Tom bluffar .
Tom fuskar .
Tom är gladlynt .
Tom är glad av sig .
Tom är munter .
Tom är förvirrad .
Tom drömmer .
Tom drunknar .
Tom är orädd .
Tom är oförskräckt .
Tom är färdig .
Tom är klar .
Tom är vänlig .
Tom sörjer .
Tom är oförarglig .
Tom är ofarlig .
Tom är hemlös .
Tom har hemlängtan .
Tom skrattar .
Tom är inte här .
Tom målar .
Tom har sagt upp sig .
Tom har kommit tillbaka .
Tom simmar .
det är Tom som bestämmer .
Höj volymen på teven .
tvätta ditt ansikte .
vi kan göra det där .
vi kan inte göra det .
vi drack en hel del .
vi drack mycket .
vi bråkar ofta .
vi kysstes bara .
vi tummade på det .
vi tog varandra i handen på det .
vi blev rånade .
vi kommer att vara där .
vi flyr .
vi är färdiga .
vi är inte säkra .
vi har slutsålt .
vi har sett henne .
var du lycklig ?
var ni lyckliga ?
vilken stor katt !
vilken stor hund !
vilket land !
så varmt det är idag !
vad varmt det är idag !
vad är de där ?
vad kan jag använda ?
vad kan det vara ?
vad kan vi göra ?
vad är det för dag ?
vilken dag är det ?
vad vann jag ?
vad bryr jag mig om det ?
vad behöver jag ?
hur är den ?
Hurdan är den ?
hur ser den ut ?
hur är det ?
hur känns det ?
var är de ?
var ligger Paris ?
var var du någonstans ?
var är min bil ?
var är mitt te ?
vem förstörde denna ?
vem förstörde det här ?
vem bor här ?
vem skulle bry sig ?
vem håller utkik ?
vem är på vakt ?
vem går på vakt ?
vem talar ?
vem pratar ?
vem är den här killen ?
vem ska man lägga skulden på ?
vem ska ges skulden ?
vems är de ?
varför frågar du ?
varför ljuger du ?
varför ljuger ni ?
ni dödade Tom .
du måste göra det .
ni måste göra det .
du verkar glad .
ni verkar glada .
ni verkar lyckliga .
du borde äta .
du kommer att klara dig .
du är inbjuden .
du är min hjälte .
du är uppriktig .
du är ärlig .
ni är uppriktiga .
ni är ärliga .
du har förändrats .
ni har förändrats .
är jag ensam här ?
tråkar jag ut dig ?
har jag någonsin fel ?
är jag i trubbel ?
är mina öron röda ?
är vi alla här ?
är vi säkra nu ?
är vi säkra än ?
är vi trygga än ?
är ni färdiga ?
är du på jobb ?
är du på jobbet ?
är du säker ?
är du avundsjuk ?
är ni avundsjuka ?
är ni avundsjuk ?
skämtar du ?
tittar du ?
är du allvarlig ?
menar du allvar ?
är du törstig ?
uppför dig .
hämta hit min väska .
ring polisen !
har jag råd med den ?
får jag vara ärlig ?
kan jag få en hund ?
får jag ta den här ?
kan jag beställa nu ?
kan jag beställa en ?
får jag parkera här ?
får jag sitta här ?
kan jag sitta här ?
kan jag lita på Tom ?
får jag prova den ?
kan jag arbeta här ?
kan Tom hjälpa oss ?
kan någon hjälpa till ?
kan den repareras ?
går den att laga ?
kan de se oss ?
kan vi äta det här ?
kan vi laga den här ?
kan vi bevisa det ?
kan vi rädda Tom ?
kan vi sitta här ?
kan vi använda den här ?
kan du känna det ?
kan du hämta Tom ?
kan du höra mig ?
hinner du ?
kan du flytta den ?
kan du läsa det ?
ser du vad det står ?
kan du hoppa över mig ?
kan du skjutsa mig ?
städa ditt rum .
stäng din bok .
stäng er bok .
stäng igen din bok .
blunda .
kom och ta mig .
kom och hälsa på oss .
kom in här .
kom in , Tom .
kom upp , Tom .
kom och prata med mig .
kom , sätt dig bredvid mig .
får jag fråga varför ?
kan jag få den ?
Kråkor är svarta .
sluta , Tom .
missade jag mycket ?
gjorde Tom det här ?
såg Tom okej ut ?
sa Tom vem ?
sa Tom varför ?
sade Tom varför ?
sa Tom ja ?
tyckte hon om den ?
köpte de den ?
gjorde du det ?
gjorde du det här ?
var det du som gjorde det här ?
hörde du det ?
tyckte du om det ?
tyckte ni om det ?
saknade du mig ?
tryckte du på den ?
läste du den ?
läste du det ?
såg du Tom ?
skrev du under det ?
skrev du på det ?
Stämde du Tom ?
tog du den ?
jag bjuder på middag .
ser jag trött ut ?
använder du droger ?
tvivlar du på mig ?
tycker ni om det ?
känns det inte bra ?
känner du dig gammal ?
känner du Tom ?
känner du till Tom ?
känner du henne ?
känner du honom ?
vet du hur ?
gillar du Tom ?
tycker du om Tom ?
älskar du Tom ?
älskar ni Tom ?
älskar du henne ?
saknar du Tom ?
saknar ni Tom ?
ser du dem ?
ser du den här ?
litar du på mig ?
Irriterar det dig ?
ser den okej ut ?
kör försiktigt .
Smaklig måltid .
alla applåderar .
alla vet .
alla är överens .
alla gjorde det .
alla bad .
alla såg det .
alla såg den .
alla är döda .
alla är här .
alla är sjuka .
följ den bilen .
Skärp dig , Tom .
skaffa ett liv , Tom .
gå in i båten .
sätt dig i båten .
Försvinn från min gräsmatta !
Åk ut ur stan .
få bort dem .
Röj undan dem .
hämta kaptenen .
hämta din mamma .
slå Tom en signal .
ge Tom ett handtag .
ge mig en munk .
ge mig någonting att dricka .
ge mig eld .
ge mig en sked .
ge mig en timme .
ge mig min käpp .
ge dem pengar .
gå ut tillbaka .
Återgå till arbetet .
gå och gör någonting .
gå och hämta din bil .
gå in i labbet .
gå och gör popcorn .
gå till läkaren .
gå till jobbet , Tom .
gå till din plats .
håll i dem .
har Tom kommit ?
har han kommit än ?
ha en bra dag .
ha en bra dag .
han började gråta .
han gjorde sin plikt .
han drack en öl .
han hade inga pengar .
han har en Toyota .
han har gått ut .
han har tio kossor .
han har tio kor .
han är en slug räv .
han är lärare .
han är ogift .
han är välavlönad .
han gillar att springa .
han ser stark ut .
han blev av med sitt jobb .
han älskar fotboll .
han älskar tåg .
han kan vara där .
han nämnde det .
han läser arabiska .
han säljer radioapparater .
han blir lätt trött .
han skriver böcker .
han håller på att bli skallig .
snälla hjälp mig .
hennes bok är röd .
hennes hår är torrt .
här är jag igen .
här är bilen .
här , prova den .
hör ni , jag kan hjälpa till .
Hallå , kan jag hjälpa till ?
hans namn är Tom .
han heter Tom .
Hissa seglen !
håll Tom åt mig .
kan du inte ge en kram ?
kan jag få en kram ?
hur mår du nu ?
hur kan vi stå till tjänst ?
hur agerade Tom ?
hur ska vi börja ?
hur smakar maten ?
hur är det med din pappa ?
hur gammal är du ?
hur gammal är den där ?
hur gammal är den här ?
hur rik är Tom ?
hur sjuk är Tom ?
hur ska det sluta ?
hur är det med Tom ?
hur går det för Tom ?
hur går det ?
jag avskyr spindlar .
det värker i hela kroppen .
jag har ont överallt .
jag gjorde det nästan .
jag är från Egypten .
jag frågade efter Tom .
det där måste ha gjort ont .
jag köpte en bok .
jag kom trea .
jag kom med Tom .
jag kan vara ärlig .
jag kan göra det nu .
jag kan köra dig .
jag kan känna det .
jag kan få in oss .
jag kan simma bra .
jag kan lita på Tom .
jag kan gå hem .
jag kan jobba sent .
jag kan inte vara säker .
jag kan inte delta .
jag kan inte tävla .
jag kan inte ställa upp .
jag kan inte göra detta .
jag kan inte låtsas .
jag kan inte bluffa det .
jag kan inte fejka det .
jag kan inte hitta den .
jag kan inte hitta det .
jag hinner inte .
jag kan inte göra det ogjort .
jag fångade en fisk !
jag lagade kvällsmat .
jag lagade middag .
jag skulle kunna göra det .
jag skulle behöva en .
jag tar gärna en .
jag gråter varje dag .
jag gjorde det en gång .
det stör mig inte .
jag körde bilen .
jag tycker om att jobba .
jag avfyrade ett skott .
jag glömde min väska .
jag hittade min bok .
jag fick en rutten en .
jag fick en som var rutten .
jag fick rabatt .
jag kom över det .
jag köpte de här åt dig .
jag fick din lapp .
jag hade min chans .
jag hade mina dubier .
jag hade mina order .
jag var tvungen att ge upp .
jag fick säga upp mig .
jag var tvungen att säga upp mig .
jag hatar min röst .
jag hatar politik .
jag hatar regn .
jag har familj .
jag har en familj .
jag har en minut .
jag har en teori .
jag har ett äpple .
jag har bevis .
jag har en till .
jag måste hålla med .
jag måste sova .
jag har två bilar .
jag har två jobb .
jag har din nyckel .
jag hörde ett brak .
jag hörde ett ljud .
jag hörde ett oljud .
jag hörde ett ljud .
jag hoppas att det regnar .
jag hoppas att den fungerar .
jag gjorde illa armbågen .
jag tänker försöka .
jag hittade den precis .
jag hittade det just .
jag hittade den just .
jag hittade det precis .
jag har just fått den .
jag har just lämnat Tom .
jag har nyligen flyttat in .
jag har just berättat det för honom .
jag kände till risken .
jag visste för mycket .
jag kan allt det här .
jag vet allt det här .
jag kan allt detta .
jag vet allt detta .
jag vet att det gör ont .
jag kan sången .
jag kan låten .
jag känner till sången .
jag känner till låten .
jag ljög om det .
jag gillar tecknat .
jag tycker om barn .
jag tycker om att klättra .
jag tycker om klättring .
jag gillar att simma .
jag tycker om att simma .
jag tycker om simning .
jag tycker om det jobbet .
jag gillar den där slipsen .
jag gillar den här koppen .
jag gillar den här hunden .
jag tycker om den här hunden .
jag tycker om att dansa .
jag tycker om dig också .
jag gillar din hund .
jag tycker om din hund .
jag gillar din hatt .
jag tycker om din hatt .
jag tände tändstickan .
jag bor i Japan .
jag bor med Tom .
jag bodde i Rom .
jag älskar barn .
jag älskar den här bilen .
jag älskar det här jobbet .
jag älskar detta jobb .
jag älskar detta arbete .
jag älskar det här arbetet .
jag älskar att skrinna .
jag älskar att undervisa .
jag älskar er båda .
jag tycker jättemycket om din väska .
din väska är jättefin .
du har jättefin hatt .
jag gjorde den där .
jag tänkte ringa .
jag träffade Tom idag .
jag träffade henne igen .
jag saknar allt det här .
jag saknar dig , Tom .
jag saknar dig också .
jag missförstod .
jag måste vara full .
jag måste vara där .
jag måste ta reda på det .
jag måste få reda på det .
jag måste hjälpa honom .
jag måste träffa Tom .
jag måste tala om det för Tom .
jag måste säga det till Tom .
jag måste berätta det för Tom .
jag behöver internet .
jag behöver en advokat .
jag behöver en minut .
jag behöver ett vapen .
jag behöver bevis .
jag behöver hans namn .
jag behöver mina tabletter .
jag behöver en till .
jag behöver lite frisk luft .
jag behöver någon .
jag behöver nycklarna .
jag behöver bandet .
jag behöver dig här .
jag behöver din bil .
jag ger aldrig upp .
jag slog aldrig Tom .
jag träffade aldrig Tom .
jag såg dig aldrig .
jag såg aldrig dig .
jag såg aldrig er .
jag såg er aldrig .
jag ser honom ofta .
jag träffar honom ofta .
jag betalade mina räkningar .
jag betalade mina skatter .
jag spelade tennis .
jag ringde i klockan .
jag läste ett brev .
jag läser ett brev .
jag litade på Tom .
jag springer varje dag .
jag joggar varje dag .
lägg av , sa jag !
jag sa det jag ville säga .
sätt dig , sa jag .
jag sa för mycket .
jag såg Tom igen .
jag såg Tom rodna .
jag såg Tom le .
jag såg Tom i dag .
jag träffade Tom i dag .
jag såg honom där .
jag såg ett idag .
jag såg den där också .
jag såg bråket .
jag såg grälet .
jag såg dig där .
jag ser ett mönster .
jag ser honom ofta .
jag ser krönet .
jag ser toppen .
jag skickade iväg Tom .
jag skickade hem Tom .
jag sov hela dagen .
jag talar svenska .
jag pratar svenska .
jag gör det fortfarande .
jag läser spanska .
jag studerar spanska .
jag pratade med Tom .
jag talade med Tom .
jag är benägen att hålla med .
jag sa det till Tom .
jag litar på er alla .
jag litar på er allihopa .
jag stängde av den .
jag vill ha en Toyota .
jag vill ha en gitarr .
jag vill ha en advokat .
jag vill ha en papegoja .
jag vill ha pengarna tillbaka .
jag vill ha ett äpple .
jag vill ha den väskan .
jag vill ha den där bilen .
jag vill ha den här väskan .
jag vill dansa .
jag föddes här .
jag var äcklad .
jag var förfärad .
jag var i Boston .
jag var ansvarig .
jag höll i trådarna .
jag var väldigt upptagen .
jag ska hjälpa dig .
jag önskar dig lycka till .
jag önskar dig lycka .
jag önskar dig allt väl .
jag önskar dig lycka till .
jag jobbar här nu .
jag jobbar här numera .
jag ska göra mitt bästa .
jag hämtar min bil .
jag går och frågar Tom .
jag kommer att gå och fråga Tom .
jag går och hämtar Tom .
jag betalar det dubbla .
jag är glad att vi träffades .
jag blir galen .
jag hjälper dig .
jag är vänsterhänt .
jag är fyndig .
jag är påhittig .
jag är rådig .
jag är fortfarande arg .
jag är trött på TV .
jag är din advokat .
jag måste iväg .
jag måste kila .
jag måste försöka .
är Tom medlem ?
är Tom så dålig ?
är Tom så usel ?
är Tom din son ?
är Tom er son ?
är någon hemma ?
andas han ?
är den giftig ?
är det giftigt ?
är hon japansk ?
är hon japanska ?
är det hälsosamt ?
är det där hälsosamt ?
är det här en radio ?
är det här korrekt ?
är det här riktigt ?
är det här etiskt ?
är det här allvarligt ?
är det måndag idag ?
det skulle kunna vara kul .
det skulle kunna vara roligt .
det måste vara jag .
den såg billig ut .
det såg billigt ut .
det såg roligt ut .
det var väldigt varmt .
det var värt det .
det är kallt i dag .
det är influensasäsong .
det är lunchdags .
det är inget problem .
det är inga problem .
det är inte en lek .
det är inte så illa .
den är utomordentlig .
det är dags att åka .
det är dags att gå .
Jesus älskar dig .
låt mig se det där .
låt mig berätta för Tom .
vi stannar här .
livet är inte lätt .
livet är inte lätt .
se dig omkring .
titta på katten .
titta bakom dig .
jag kanske stannar .
Blanda Tom en drink .
min hund sprang iväg .
min hund har sprungit iväg .
jag har ont i halsen .
ingen blev sjuk .
ingen är där .
ingen skadades .
ingenting är gratis .
gå och lägg dig nu .
gå och lägg er nu .
öppna flaskan .
öppna munnen !
öppna munnen .
Varsågod och sitt ner .
Läs detta först .
Läs det här först .
regler är regler .
spara en munk till mig .
säg nej till droger .
hajar äter fisk .
hon hade en radio .
hon bor ensam .
hon tittade bort .
hon gick ut .
hon väckte honom .
sitt rakt .
så vad ska jag göra ?
våren är här .
Våran har kommit .
våren är kommen .
berätta en historia .
berätta en saga .
säg vem som vann .
den bilen är hans .
det där är ett hjärta .
det där är ett bord .
det där är hans bil .
det där är en pagoda .
det är gammal skåpmat .
luften är fuktig .
svaret är nej .
bilen är blå .
hunden är död .
det finns ingen tvål .
de är skådespelare .
de dog unga .
de gick tidigt .
de bor där .
de förlorade igen .
de blev tokiga .
den här bilen är hans .
det här är min öl .
det här är mitt öl .
det här är mitt skepp .
detta är min fru .
det här är slutet .
kasta den till Tom .
att fela är mänskligt .
Tom hade inget emot det .
Tom överdrev .
Tom klädde på sig .
Tom förlovade sig .
Tom blev ivrig .
Tom hade ingenting .
Tom har anlänt .
Tom har kommit .
Tom har förändrats .
Tom har rymt .
Tom har kaniner .
Tom hatade att ljuga .
Tom hatar lögnare .
Tom hatar lögnhalsar .
Tom hatar opera .
Tom är en hippie .
Tom är bedårande .
Tom är förtjusande .
Tom är upprörd .
Tom är irriterande .
Tom är konstnärlig .
Tom är atletisk .
Tom har autism .
Tom är autistisk .
Tom bluffar .
Tom är charmig .
Tom är kreativ .
Tom är trovärdig .
Tom är kultiverad .
Tom är finkänslig .
Tom är sinnessjuk .
Tom är vansinnig .
Tom är flitig .
Tom är illojal .
Tom är skild .
Tom är villrådig .
Tom är dyblöt .
Tom är genomvåt .
Tom är orädd .
Tom är vänlig .
Tom skrattar .
Tom är inte här .
Tom målar .
Tom är fortfarande uppe .
Tom är fortfarande vaken .
Tom simmar .
det är Tom som bestämmer .
Tom är chef .
Tom är för långsam .
Tom är på övervåningen .
Tom har det bra ställt .
Tom är inte petig .
Tom är inte glad .
Tom är inte småaktig .
Tom dödade Mary .
Tom lämnade ett meddelande .
Tom ljög för dig .
Tom såg bra ut .
Tom ser arg ut .
Tom ser glad ut .
Tom ser trött ut .
Tom saknar Mary .
Tom verkade borta .
Tom verkade vilse .
Tom verkade trevlig .
Tom verkar uttråkad .
Tom stannade hemma .
Tom berättade ett skämt .
Tom berättade en vits .
Tom bleknade .
Tom blev blek .
Tom var tillgiven .
Tom var som jag .
Tom var min hjälte .
Tom flämtade .
Tom flåsade .
Tom stönade .
Tom hade helt rätt .
Tom är genialisk .
Tom är bekymrad .
Tom är vid medvetande .
Tom är vid sans .
Tom är övertygad .
Tom är farlig .
Tom är desperat .
Tom är annorlunda .
Tom är imponerad .
vänta en sekund .
tvätta händerna .
se upp var du går .
vi är i Paris .
vi är studenter .
vi tittar .
vi måste flytta .
vi måste förflytta oss .
vi älskar picknickar .
vi måste hitta den .
vi måste hitta det .
vi borde studera .
vi var oroliga .
vi jobbar för Tom .
vi är anpassningsbara .
vi kan anpassa oss .
vi är flexibla .
vi är annorlunda .
vi är olika .
vad kan Tom göra ?
vad gjorde Tom ?
vad sa han ?
vad sade han ?
vad fick vi ?
vad gör de ?
vad har vi ?
vad vet vi ?
hur är han ?
Hurdan är han ?
vad är det , Tom ?
vad saknas ?
vad dödade Tom ?
vad var det som Tom dödade ?
vad skrämde dig ?
vad fanns inuti ?
vad heter han ?
vad finns där inne ?
vad finns på insidan ?
vad handlar det om ?
vad är min belöning ?
vad är det som är så kul ?
vad är det som är så roligt ?
vad är klockan ?
vad är den här till ?
vad används den här till ?
vad har du ?
när kan vi äta ?
när ska vi gå ?
vart gick han ?
var är väskan ?
vem är den killen ?
vem är den där killen ?
vem är den där mannen ?
vem tog emot det ?
du vart lurad .
du ser dum ut .
ni borde stanna .
du skrämde mig .
du kommer snart att dö .
ni är bedårande .
du är förtjusande .
ni är förtjusande .
du är en idiot .
du är arrogant .
ni är arroganta .
du är atletisk .
ni är atletiska .
du babblar .
du pladdrar .
du är oartig .
ni är oartiga .
du är mitt barn .
du kör så mycket med folk .
du domderar så mycket .
du är så kinkig .
du är så kräsen .
du kommer med undanflykter .
du är begåvad .
din katt är tjock .
er katt är tjock .
en taxi står och väntar .
en hund skäller .
en tjej ringde mig .
får jag sparken ?
vem som helst kan göra det .
är de förälskade i varandra ?
är de där till mig ?
är de där för mig ?
är de där åt mig ?
är vi färdiga här ?
ska vi åka långt ?
ska vi gå långt ?
är du amerikan ?
är du japansk ?
är du golfspelare ?
är du förälder ?
är du präst ?
är du en idiot ?
Rodnar du ?
går det bra för dig ?
tänker du gå in ?
är du i Paris ?
är ni i Paris ?
är du min fiende ?
är du ny här ?
är du ombord ?
använder du droger ?
har ni öppet nu ?
sover du ?
har du för kallt ?
har du för varmt ?
är ni två upptagna ?
är du där uppe ?
kom dit vid tolv .
hämta in den , Tom .
kom igen , Tom .
hämta min käpp .
hämta hit dem .
borsta tänderna .
borsta dina tänder .
borsta era tänder .
kan jag vara till hjälp ?
kan jag få en öl ?
får jag stiga upp nu ?
får jag gå och surfa ?
kan jag få en kram ?
kan jag få tre ?
kan jag lita på dem ?
kan Tom gå först ?
går detta att utföra ?
kan detta vara sant ?
kan vi ta med Tom ?
får vi också komma ?
kan vi hjälpa dem ?
kan vi gå nu ?
kan vi bo här ?
kan vi prata här ?
kan vi lita på dig ?
kan du fånga mig ?
kan du ta reda på det ?
kan du bevisa det ?
kan du rädda Tom ?
kan du se det där ?
kan du se dem ?
kan ni se dem ?
kan du tala högre ?
kan du stoppa Tom ?
kan du inte se det ?
kan du inte se den ?
städa upp det , Tom .
klättra upp till toppen .
kom och hjälp oss .
kom igen , rör på påkarna .
kom ut med oss .
kom och spring med mig .
Fortsätt gräva .
Fortsätt arbeta .
Behärska dig .
kan det vara sant ?
bjöd jag in dig ?
skrev jag det där ?
bet Tom dig ?
blev Tom skadad ?
skadades Tom ?
slog Tom Mary ?
betalade Tom också ?
Knuffade Tom dig ?
Pressade Tom dig ?
har Tom sänt dig ?
hittade de den ?
hade de den ?
sa de hur ?
sade de hur ?
sa de varför ?
sade de varför ?
tog du med den ?
hittade du Tom ?
gick du vilse ?
fick du det ?
förstod du det där ?
hade du roligt ?
hade du kul ?
dödade du Tom ?
kände du Tom ?
träffade du honom ?
svimmade du ?
sov du bra ?
berättade du för Tom ?
varnade du Tom ?
får jag ett pris ?
ser jag normal ut ?
ser jag dum ut ?
ser jag ut som trettio ?
är det bacon jag känner lukten av ?
gör som du vill .
gör det igen , Tom .
gör det en gång till .
gör vad du vill .
gör vad du vill .
klandrar du Tom ?
Förebrår du Tom ?
lägger du skulden på Tom ?
Hänger du med på vad jag menar ?
har du dem ?
känner du dem ?
gillar du golf ?
gillar du snö ?
tycker du om snö ?
gillar du dem ?
tycker du om vin ?
bor du här ?
bor ni här ?
menar du det ?
behöver du dem ?
spelar du golf ?
läser du på läppar ?
säljer ni vin ?
litar du på Tom ?
vill du ha fisk ?
vill du ha barn ?
vill du ha mera ?
vill du ha litet ?
vill du ha dem ?
är du anställd här ?
är det Tom som har den ?
tycker Tom om mig ?
var inte så lat .
drick inte det där .
Överdriv inte .
inte så fort !
ingen orsak .
prata inte med mig .
tala inte med mig .
rita en linje här .
ät dina grönsaker .
alla jämrar sig .
alla skrattar .
alla log .
alla stannade .
alla väntade .
alla är upptagna .
alla flydde .
alla ska gå .
alla är tysta .
alla är där .
slåss som en man !
Tanka full tank .
glöm henne .
kom in och kör .
sätt dig i lastbilen .
hämta lite vin åt mig .
ta lite åt mig också .
gå bort från min veranda .
gå ner på golvet .
sätt igång och jobba , Tom .
ge Tom någonting att dricka .
ge Tom pistolen .
ge det en chans .
ge den en minut .
ropa på mig .
vänta en stund .
ge mig ett ögonblick .
ge mig mina pengar .
ge mig en timme .
ge mig en till .
ge mig den där pistolen .
ge mig det där geväret .
ge mig den där nyckeln .
ge mig filen .
ge mig vinet .
ge mig den här hatten .
ge mig din arm .
ge det här till Tom .
ge oss en chans .
ge oss ett ögonblick .
ge oss en sekund .
säg det bara .
säg det nu .
gå raka vägen hem .
gå och lägg dig , Tom .
gå till garaget .
ta ett paraply .
ta en åt mig också .
ge mig en servett .
har Tom blivit matad ?
är det någon som har dött ?
få Tom att ringa mig .
ha ett bra liv .
ha en jättebra dag .
ha en fantastisk dag .
ha ett bra liv .
ha ett trevligt liv .
ha en trevlig simtur .
har du träffat Tom ?
har ni beställt ?
har du läst den ?
har ni två träffats ?
hon började springa .
han bar sig illa åt .
han bröt armen .
han föll baklänges .
han hittade min cykel .
han hade få tänder .
han är italienare .
han är akrobat .
han har problem .
han tycker om djur .
han tycker om att sjunga .
han tycker om att simma .
han tycker om djur .
han gav inget svar .
han måste älska dig .
han spelade tennis .
han såg hennes video .
han blir rädd lätt .
han blir lätt rädd .
han sov hela dagen .
han talar arabiska .
han talar franska .
han tog sin tid .
han vill ha en iPad .
han var i Frankrike .
han var fängslad .
han har glasögon .
han har på sig glasögon .
han jobbar söndagar .
han är en gentleman .
han är vid hennes sida .
han är din vän .
han är din kompis .
här , prova min penna .
här , använd min penna .
Hallå , är det du som är Tom ?
Hallå där , vem är du ?
vänta ett ögonblick .
vänta lite nu .
håll det där åt mig .
kan jag få en puss ?
hur smakar äggen ?
hur mår du ?
hur går det för dig ?
hur mår ni ?
hur kommer det sig att du frågar ?
hur kunde Tom veta om det ?
hur såg Tom ut ?
hur dog de ?
hur visste du ?
hur ska jag göra det ?
hur ska jag göra det här ?
hur ska jag svara ?
hur känner de sig ?
hur kan de veta det ?
hur ser de ut ?
hur ser det ut ?
hur fungerar det ?
så pinsamt !
hur kan det här vara rättvist ?
hur stor var den ?
hur mycket är det där ?
hur var det idag ?
hur var föreställningen ?
hur var resan ?
hur var din tupplur ?
vad du har växt !
jag håller med Tom .
jag gjorde det redan .
jag tycker också om katter .
jag gör alltid sådär .
jag kommer ifrån Ryssland .
jag kommer från Ryssland .
jag är ifrån Ryssland .
jag är ingen häxa .
jag började gripas av panik .
jag börjar imorgon .
jag slår vad om att Tom har glömt .
jag slår vad om att det var Tom .
det är jag som bestämmer .
jag kom tillbaka hem .
jag kom för att säga hej .
jag kan vara tålmodig .
jag kan bära den där .
jag kan också göra det .
jag kan få in dig .
jag kan ta hand om Tom .
jag kan nämna några namn .
jag kan känna lukten av rädsla .
jag kan inte röra det ur fläcken .
jag kan inte flytta på det .
jag bryr mig om Tom .
jag skulle kunna hjälpa Tom .
jag skulle kunna hjälpa dig .
jag skulle kunna döda dig .
jag skulle kunna kyssa dig .
jag kunde inte sova .
jag kunde inte stå .
jag gjorde det för Tom .
jag gör mitt jobb väl .
jag känner inte Tom .
jag känner inte honom .
jag kör en hybrid .
jag kör en hybridbil .
jag blev underkänd i provet .
jag känner mig självsäker .
jag mår ganska dåligt .
jag känner mig så vacker .
jag känner mig så dum .
jag känner mig väldigt kall .
jag kände mig skräckslagen .
jag fyllde koppen .
jag fyllde på i koppen .
jag glömde kartan .
jag hittade mina skor .
jag fann mina skor .
jag hittade nycklarna .
jag hittade den här .
jag gav det ett försök .
jag sa upp mig .
jag fattar vad du menar .
jag fick en bra en .
jag kom hem först .
jag skaffade en åt oss .
jag blev betalad i dag .
jag har haft en tung dag .
det har varit en tung dag .
jag hade huvudvärk .
vi var tvungna att göra det .
jag var tvungen att gå hem .
jag hatar kemi .
jag hatar min familj .
jag hatar min syster .
jag hatar överraskningar .
jag hatar den idén .
jag hatar det här spelet .
jag hatar den här sången .
jag hatar den här låten .
jag avskyr dig som pesten .
jag har en kommentar .
jag har ett diplom .
jag har en akademisk examen .
jag har en brödrost .
jag har en husvagn .
jag har varit upptagen .
jag har blå ögon .
jag har blåa ögon .
jag har god hörsel .
jag har god syn .
jag har goda nyheter .
jag har juryplikt .
jag har mina begränsningar .
jag har mina order .
jag har mina saker .
jag måste avbryta .
jag måste ändra på mig .
jag måste gå nu .
jag måste bege mig nu .
jag måste ge mig av nu .
jag måste gå ut .
jag måste prova det .
jag har din fil .
jag hörde det på tv .
jag hörde klockan .
jag hoppas att jag överlever .
jag hoppas att Tom är okej .
det insisterar jag på .
jag har alldeles nyss gett Tom sparken .
jag har alldeles nyss avskedat Tom .
jag fick precis sparken .
jag öppnade den precis .
jag för dagbok .
jag för en journal .
jag höll mig för mig själv .
jag kände till riskerna .
jag vet att jag har fel .
jag känner till den där blicken .
så mycket vet jag .
det där vet jag .
jag känner till det namnet .
jag vet det , Tom .
jag kan rutinen .
jag vet hur det går till .
jag känner ägaren .
jag vet vad det rör sig om .
jag vet att du försökte .
jag känner igen ditt ansikte .
jag åkte för tidigt .
jag tycker om choklad .
jag tycker om hundar också .
jag gillar grönt te .
jag tycker om grönt te .
jag tycker om att resa .
jag gillar ditt hår .
jag bor i lägenheten bredvid .
jag älskar astronomi .
jag älskar min mamma .
jag älskar den sången .
jag älskar den här delen .
jag älskar denna del .
jag älskar den här staden .
jag älskar denna stad .
jag älskar att resa .
jag älskar dina ögon .
jag älskar ditt hår .
jag älskade pjäsen .
jag älskade dig en gång .
jag gjorde en snögubbe .
jag gjorde frukost .
jag gör upp reglerna .
jag får dig att le .
jag kan bli vald .
jag kanske inte återvänder .
jag mjölkade kon .
jag måste bege mig nu .
jag måste ge mig av nu .
jag måste lämna dig .
jag behöver Tom levande .
jag behöver en ny .
jag behöver en röd penna .
jag behöver hela rubbet .
jag behöver ett svar .
jag behöver frisk luft .
jag behöver mer hjälp .
jag behöver mer tid .
jag behöver det där bandet .
jag behöver sanningen .
jag måste se den .
jag måste varva ner .
jag tyckte aldrig om den .
jag tar aldrig sovmorgon .
jag äter ofta här .
jag behöver bara hälften .
jag äger den här affären .
jag har planterat ett träd .
jag föredrar att gå .
jag läste etiketten .
jag menar det verkligen .
jag saknar det verkligen .
jag vägrar hjälpa till .
jag vägrar hjälpa .
jag vägrar arbeta .
Strunta i det , sa jag .
bry dig inte om det , sa jag .
stanna här , sa jag .
gå undan , sa jag .
stig åt sidan , sa jag .
jag såg när Tom kom .
jag såg lite rök .
jag var hos läkaren .
jag såg dig gråta .
jag sköt hästen .
jag borde stämma Tom .
jag talade inför klassen .
jag tycker fortfarande om Tom .
jag tycker fortfarande om dig .
jag saknar Tom fortfarande .
jag tror att Tom gick .
jag tog pengarna .
jag tog fotot .
det tvivlar jag verkligen på .
jag hoppas verkligen inte det .
jag vill ha en tvättbjörn .
jag vill ha en sparkcykel .
jag vill ha mera mat .
jag vill resa .
jag var en främling .
jag hade bara tur .
jag var ganska upptagen .
jag var så nervös .
jag var väldigt glad .
jag var mycket glad .
jag tvättade bilen .
jag kommer inte att vara tyst .
jag kommer inte att behöva dig .
jag kommer inte att behöva er .
jag arbetade för Tom .
jag skulle inte göra det .
det är nog bäst att jag går .
jag hade sagt nej .
jag skulle vilja hjälpa till .
jag är hos Tom .
jag kommer att straffas .
jag ska kolla igen .
jag kommer att få tillbaka den .
jag ska hämta min jacka .
jag ska ta min jacka .
jag ska hämta min rock .
jag ska hämta min kappa .
jag ska ta min kappa .
jag hämtar mina nycklar .
jag hämtar nycklarna .
jag ska hämta mina nycklar .
jag ska hämta nycklarna .
jag kommer över det .
jag kommer nog över det .
jag hämtar bilen .
jag ska hämta bilen .
jag går och hämtar lite .
jag går och hämtar det .
jag går in först .
jag ska gå och handla .
jag ska gå och shoppa .
jag går den här vägen .
jag ska gå med Tom .
jag följer med dig .
jag kommer att följa med dig .
jag ska följa med dig .
jag tar hand om det här .
jag kommer att ta hand om det här .
jag ska ta hand om det här .
jag hämtar upp Tom .
jag kommer att hämta upp Tom .
jag ska hämta upp Tom .
jag pratar med Tom .
jag ska prata med Tom .
jag kommer att prata med Tom .
jag ska göra mitt bästa .
jag ska vänta en vecka .
jag är lite hungrig .
jag är redan rik .
jag är upptagen i kväll .
det är roligt att kunna hjälpa till .
jag ska försöka .
jag kommer att försöka .
jag är på vinden .
jag är på vindsvåningen .
jag är ingen tiggare .
jag är inte läkare .
jag är inte så trött .
jag är på din sida .
jag är stolt över dig .
jag är också pensionerad .
jag är trött på det här .
jag har fått nog av det här .
jag är liksom upptagen .
jag stannar här .
jag är väldigt törstig .
jag är din bror .
jag är er bror .
jag har sällskap .
jag måste få veta .
jag måste sluta .
jag måste stanna .
jag har tappat bort min penna .
jag har aldrig röstat .
är Tom säker ?
är Tom där ute ?
är Tom där än ?
smittar det ?
är det för svårt ?
det kostar två euro .
det är din rättighet .
det fick mig att skratta .
det kanske blir regn snart .
det var inte en tävling .
det får duga .
det måste duga .
det är en dålig vana .
det är allt vi har .
den är allt vi har .
den är bekväm .
det är bekvämt .
det är dimmigt i dag .
det är intressant .
det är mitt beslut .
beslutet är mitt .
den är inte till dig .
det är inte till dig .
den är inte till er .
det är inte till er .
det är inte från mig .
den är inte från mig .
det är bara en bok .
det är ganska kallt .
den är begagnad .
den är second hand .
det är värt ett försök .
gör bara som jag säger .
Posta det här brevet .
gör ditt val .
får jag öppna en burk ?
min bil är en tysk bil .
mina ögon är blå .
mina ögon är ömma .
min far är inte hemma .
min far röker .
mina fötter är ömma .
mitt glas är fullt .
min inkorg är full .
mina nycklar är borta .
det gör ont i mitt ben nu .
det gör ont i benet nu .
mitt ben är brutet .
min näsa kliar .
min tid är kommen .
ingen får avlägsna sig .
nu känner jag mig trött .
kom med mig nu .
ge tillbaka den nu .
ge mig det där nu .
ge mig den där nu .
gå in nu .
låt mig tänka nu .
se nu på der här .
skicka saltet .
snälla kör in till trottoarkanten .
rödvin , tack .
skolan är tråkig .
hon dog 1960 .
hon gillar att springa .
hon kanske inte kommer .
så vad hände ?
spindlar skrämmer mig .
stanna bilen nu !
ta hand om Tom .
säg åt Tom att vänta .
det är obotligt .
det där är min hemlighet .
det där är inte billigt .
det är irrelevant .
det är inte relaterat .
det är jättefint !
det är fantastiskt !
det var roligt att höra !
det är min bok .
hunden är döende .
hunden är smart .
Juryn är oenig .
Bucklan var min .
Pottan var min .
Krukan var min .
burken var min .
Kannan var min .
Haschet var mitt .
de bor här nära .
de bor i närheten .
de tog i hand .
de skakade hand .
de tackade Gud .
de var hjältar .
de är gräsliga .
de är förfärliga .
de är inte upptagna .
de kommer med undanflykter .
de slingrar sig .
de överstegrar .
de är likadana .
den här pojken är lat .
den här hunden är min .
det här är bevis .
det här är min häst .
detta är min häst .
det här är mitt hus .
det här är rödvin .
det här är för svårt .
det här är inte rätt .
detta är inte rätt .
detta stämmer inte .
det här stämmer inte .
det här blir kul .
Tom svarade ja .
Tom åt sig mätt .
Tom åt så mycket han orkade .
Tom studsade tillbaka .
Tom kom för att hjälpa .
Tom kan höra dig .
Tom kan höra er .
Tom kan inte vägra .
Tom kan inte neka .
Tom kan inte säga nej .
Tom klättrade ner .
Tom vet inte .
Tom förklarade det .
Tom sneglade neråt .
Tom blev arresterad .
Tom blev förvirrad .
Tom har ambitioner .
Tom har barn .
Tom har fräknar .
Tom har undantagsrätt .
Tom har immunitet .
Tom har åkt fast för rattfylleri två gånger .
Tom hatade att gå i skola .
Tom hatade skolan .
Tom avskyr oliver .
Tom hjälpte mycket .
Tom är en beatnik .
Tom är en hipster .
Tom är en stamkund .
Tom är en stamgäst .
Tom är fast anställd .
Tom är ambitiös .
Tom är föräldralös .
Tom är ett föräldralöst barn .
Tom är engagerad .
Tom är kompetent .
Tom är skicklig .
Tom är bekymrad .
Tom är säker .
Tom är nöjd .
Tom är belåten .
Tom är artig .
Tom är hövlig .
Tom är förtjust .
Tom är nedstämd .
Tom är deprimerad .
Tom är desperat .
Tom är oärlig .
Tom ligger i koma .
Tom är olycklig .
Tom är förtvivlad .
Tom är min brorson .
Tom är min systerson .
Tom är nonchalant .
Tom är för ung .
Tom är inte rädd .
Tom gillar det hett .
Tom gillar det varmt .
Tom gillar den varm .
Tom bor här nära .
Tom tittade framåt .
Tom såg bra ut .
Tom ser road ut .
Tom ser skyldig ut .
Tom slutade röka .
Tom säljer kaffe .
Tom borde vara okej .
Tom stod förstelnad .
Tom ville ha ett jobb .
Tom ville ha ett arbete .
Tom ville ha pengar .
Tom vill ha en kyss .
Tom vill ha en puss .
Tom blev kidnappad .
Tom blev bortförd .
Tom blev bortrövad .
Tom blev arresterad .
Tom försvann .
Tom kommer att hitta den .
Tom lyssnar inte .
Tom är i våningen under .
Tom är i nedre våningen .
Tom är halsstarrig .
Tom är hårdnackad .
Tom är egensinnig .
Tom är styvsint .
sänk volymen på teven .
gå långsammare .
blev Tom mördad ?
det var väl trevligt ?
vi behöver alla kärlek .
alla behöver vi kärlek .
det kan vi inte göra .
vi har inget socker .
vi måste göra det .
vi bor tillsammans .
vi måste skynda oss .
vi vill bara ha er .
vi vill endast ha dig .
vi vill endast ha er .
vi springer varje dag .
vi var så nära .
vi var så stolta .
vi var väldigt ledsna .
vi önskar er lycka till .
vi önskar dig lycka till .
vi går och hämtar Tom .
vi är lite sena .
vi är aningens sena .
vi skär ned .
vi har problem .
vi är i trubbel .
vi är illa ute .
vi är i knipa .
vi har råkat illa ut .
vi köper inte .
jag är här .
jag är precis här .
blev du beskjuten ?
vilken usel film !
vilken dålig film !
vilken söt flicka !
vilken söt tjej !
vilken usel dag !
vilken fyndig idé !
vad kan jag ta med ?
vad kan Tom säga ?
vad kan de göra ?
vad sa Tom ?
vad sade Tom ?
vad betydde det ?
vad innebar det ?
vad köpte du ?
vad träffade du ?
vad såg du ?
vad ska jag göra nu ?
vad hatar du ?
vad har du ?
vad vet du ?
vad älskar du ?
vad söker du ?
vad vill du ?
vad vill du ha ?
vad är allt det där ?
vad är allt det här ?
vad är allt detta ?
vad har vi för plan ?
vad är det här för ?
vad är det här till ?
vad är detta för ?
vad är detta till ?
hur var det ?
vad har Tom hittat ?
vad är haken ?
vad är orsaken ?
Vadan denna panik ?
vad är ditt namn ?
vad är er plan ?
vad har du gjort ?
vad har ni gjort ?
när ska ni gå ?
när ska du gå ?
vart är jag på väg ?
var är vi nu ?
vart gick Tom ?
var är alla ?
var är allihopa ?
var är allesammans ?
var är min telefon ?
var är chefen ?
var är utgången ?
var ligger utgången ?
vem vet inte ?
vem målade den där ?
vem är nummer ett ?
vem är det som är nummer ett ?
varför är du hemma ?
varför är ni hemma ?
varför slutade ni ?
varför gör du det ?
kommer det ta lång tid för dig ?
äggulor är gula .
du kan skylla på mig .
ni kan skylla på mig .
du får skylla på mig .
ni får skylla på mig .
du förtjänar det här .
du skulle bara veta .
du behöver terapi .
du verkar frånvarande .
du borde sova .
ni borde sova .
du är misslyckad .
du är farlig .
du är annorlunda .
du är väldigt söt .
du har blivit tjock .
din hund är här .
er hund är här .
du är röd i ansiktet .
en hund sprang .
det regnade hårt .
kommer jag att dö ?
finns jag på den listan ?
är jag välkommen här ?
Ammoniak är en bas .
är de galna allihopa ?
är de i Paris ?
ska vi gå hem ?
är vi illa ute ?
är du tvåspråkig ?
är du uttråkad ännu ?
är du klar , Tom ?
ska du ut ?
är du också hemma ?
är du skadad , Tom ?
är du i fara ?
lyssnar du ?
är du vår fiende ?
är du där ute ?
är du klar nu ?
är ni klara nu ?
är du färdig ännu ?
är du klar ännu ?
är det säkert att du är okej ?
är du säker , Tom ?
är du för trött ?
är inte vi vänner ?
är inte du kock ?
är inte du köksmästare ?
var ärlig mot mig .
hämta in Tom .
köp lite godis åt mig .
får jag fråga varför inte ?
får jag fråga varför ?
kan jag fråga varför ?
kan jag göra det idag ?
får jag göra det idag ?
kan jag få en puss ?
kan jag få skjuts ?
kan jag hämta dig ?
får jag träffa Tom nu ?
får jag se något ID @-@ kort ?
kan jag tala med Tom ?
kan Tom få en hund ?
kan vi komma närmare ?
kan vi börja om från början ?
har du råd med det ?
kan du svara på det ?
kan du slå det ?
kan du frysa ner den ?
kan du frysa ned den ?
kan ni frysa ned den ?
kan du höra dem ?
hör du dem ?
hör ni dem ?
kan ni höra dem ?
kan du ta bort den ?
kan du stanna länge ?
kan du ta över ?
kan du lita på Tom ?
kan du se efter Tom ?
kan vi inte berätta för Tom ?
kan vi inte säga det till Tom ?
kan du inte göra det ?
kan ni inte göra det ?
kolla in den , Tom .
julen är här .
städa upp litet .
kom och sätt dig .
kom tillbaka hit .
kom tillbaka .
kom ner hit .
kom ut därifrån .
kom och spela med oss .
kom och lek med oss .
kom och hälsa på mig igen .
kom och bo hos mig .
kan det vara Tom ?
kan du göra det ?
kan ni hjälpa oss ?
kan du hjälpa oss ?
kan du läsa det ?
kan du läsa upp det ?
coola ner , Tom .
gjorde jag allt det där ?
kom Tom tillbaka ?
kom Tom hit ?
kom Tom hem ?
gjorde Tom Mary illa ?
såg Tom upptagen ut ?
sa Tom var ?
stannade Tom länge ?
vann Tom igen ?
gjorde de dig illa ?
sa de när ?
sade de när ?
har du ritat det där ?
kände du det där ?
hörde du det där ?
kysste du Mary ?
Pussade du Mary ?
har du gjort den här ?
menade du det ?
märkte du det ?
läste du det där ?
läste du den där ?
spelade du in det ?
har du saltat det här ?
Saltade du det här ?
skickade du dem ?
sköt du Tom ?
Fotograferade du Tom ?
skrev du under det här ?
skrev du på det här ?
har du väntat länge ?
väntade du länge ?
tvättade du den där ?
förtjänar jag det här ?
har jag feber ?
behöver jag opereras ?
har de det ?
tycker de om vin ?
arbetar de här ?
håller du med , Tom ?
dricker du , Tom ?
skrattar du någonsin ?
sover du någonsin ?
röker ni ?
har du bevis ?
kan du latin ?
vet du var ?
tycker du om godis ?
tycker du om lever ?
gillar du lever ?
tycker du om opera ?
tycker du om päron ?
tycker du om de här ?
behöver du pengar ?
behöver ni pengar ?
måste du gå ?
säljer ni frukt ?
bryr du dig fortfarande ?
vill du ha ett jobb ?
vill du ha ett arbete ?
gör ditt bästa , Tom .
tycker Tom om det ?
njuter Tom av det ?
har Tom en ?
vet Tom än ?
bor han här ?
gör det väldigt ont ?
gör det dig upprörd ?
får jag inte en kram ?
var inte barnslig .
gör inte om det .
ge inte upp nu .
berätta inte för någon .
rör inte dem .
tycker du inte om mig ?
alla hurrade .
alla överlevde .
allt är gratis .
allt är här .
stanna gärna .
fyll igen diket .
hämta lite mat åt Tom .
lämna Tom i fred .
kom ut tillbaka .
gå tillbaka upp dit .
kom in fort .
sitt upp på din häst .
kom hit nu .
gör dig färdig för att gå till sängs .
vila dig lite nu .
hämta deras vapen .
ta hit deras vapen .
vakna , allesamman .
gå och klipp dig .
hämta din anteckningsbok .
ge pappa en puss .
ge Tom en chans .
ge Tom en dollar .
ge Tom en minut .
ge Tom ett ögonblick .
ge Tom en sekund .
ge Tom hans nycklar .
ge den lite tid .
ge mig lite tid .
ge mig den där käppen .
ge mig geväret .
ge mig klockan .
ge mig ditt bälte .
ge mig din hand .
hjälp oss lite .
gå och sov en stund .
gå någon annanstans .
gå hem till Tom .
gå till Toms hus .
gå och tvätta ansiktet .
håll dig till sanningen .
har Tom blivit skadad ?
har Tom skadats ?
har Tom också gått ?
har Tom sett den här ?
har Tom sett det här ?
har Tom berättat för Mary ?
har Tom sagt det till Mary ?
ta någonting att dricka , Tom .
har de gjort det ?
har de rymt ?
har du sett Tom ?
har du sett någon ?
han utpressade mig .
han fångade en mus .
han dog i fjol .
han lyssnar inte .
han kör en Lotus .
han gav henne en låda .
han hade ont i huvudet .
han är en storätare .
han är en gentleman .
han textade mig nyss .
han höll det hemligt .
han hemlighöll det .
han hemlighöll den .
han vet för mycket .
han åkte till Paris .
han bor i Kyoto .
han ser efter oss .
han ser bekant ut .
han förlorade synen .
han behöver en stege .
han erkände sig skyldig .
han erkände .
han undervisar i arabiska .
han berättade sanningen .
han sade sanningen .
han reser runt .
han vred om min arm .
han utövade påtryckningar på mig .
han var förkrossad .
han var väldigt trött .
han vann allt .
han jobbar för mycket .
han drar ifrån .
han sitter på tåget .
hennes dröm är över .
hennes hud var varm .
här är nycklarna .
här är vi igen .
var så god , Tom .
här är ett exempel .
här är mitt kvitto .
Hallå , lyssna på mig .
hör ni , se på det där .
Hallå , var är vi ?
Hallå , var är vi någonstans ?
hans historia är sann .
Älskling , jag älskar dig .
Älskling , är du okej ?
ska vi ta oss en bit mat ?
hur illa kan det vara ?
hur dåligt kan det vara ?
hur dålig kan den vara ?
hur kan jag mäta mig med det ?
hur ska det här kunna hjälpa ?
hur kommer vi in ?
hur gjorde Tom det ?
hur svarade Tom ?
hur hade Tom sovit ?
hur lät Tom ?
hur kunde de veta om det ?
hur kunde de veta det ?
hur gissade du ?
hur ska jag äta det här ?
hur ska man äta det här ?
hur kommer jag tillbaka ?
hur ska jag hjälpa Tom ?
hur ska jag stoppa Tom ?
hur klarar du det ?
hur lyckas du ?
hur kan Tom veta det ?
hur ser Tom ut ?
hur smakar det ?
hur långt for den ?
hur rik är du ?
hur speciell är den ?
hur trött är du ?
hur var festen ?
hur var dejten ?
hur var träffen ?
hur har din vecka varit ?
det är ju jättekonstigt .
hur mår din mor ?
hur mår din mamma ?
jag sköt dig nästan .
jag hittade också den här .
jag tycker också om godis .
jag är en hundmänniska .
jag är vegetarian .
jag är alldeles förvirrad .
jag är redan sen .
jag äter frukt .
jag är inte så glad .
jag uppskattar det .
jag åt en hamburgare .
jag tror på kärleken .
du är säkert upptagen .
jag slår vad om att du är upptagen .
jag köpte en kaktus .
jag krossade hans hjärta .
jag har byggt den själv .
jag stötte på Tom .
jag kom tillbaka tidigt .
jag kom från Kina .
jag kan acceptera det .
det kan jag acceptera .
det kan jag svara på .
jag kan svara på det .
jag kan knappt röra mig .
jag kan räkna .
jag kan åka med tåg .
jag kan ta hand om det där .
jag kan slå ett samtal .
jag kan betala i förskott .
jag kan skydda dig .
jag kan cykla .
jag kan klara upp det här .
jag känner lukten av rök .
det luktar rök .
jag kan fortfarande strida .
jag kan fortfarande slåss .
jag kan fortfarande kämpa .
jag kan bekräfta det där .
det kan jag bekräfta .
jag kan inte förneka det .
jag kan inte göra det nu .
jag kan inte behålla det här .
jag kan inte behålla den här .
jag kan inte lämna dig .
jag bryr mig om det .
jag bryr mig om det här .
det här betyder mycket för mig .
jag brydde mig om Tom .
jag chartrade ett jetplan .
jag checkade in mina väskor .
jag städade mitt rum .
jag stängde porten .
jag skulle kunna sälja den här .
jag skulle kunna vara din handledare .
jag kunde inte säga nej .
jag gjorde Tom en tjänst .
jag gjorde mycket idag .
jag gjorde det här själv .
jag dödade inte Tom .
jag klandrar dig inte .
jag känner mig inte sjuk .
jag tycker inte om hundar .
jag tycker inte om ägg .
jag gillar inte ägg .
jag tycker inte om det .
jag tycker inte om det där .
jag gillar det inte .
jag behöver ingen hjälp .
jag behöver dem inte .
jag har inget behov av dem .
jag litar inte på dig .
jag vill inte ha det här .
jag vill inte ha den här .
jag vill inte ha denna .
jag vill inte ha detta .
jag kör en Porsche .
jag har jättedåligt samvete .
jag känner mig sårbar .
jag glömde min handväska .
jag hittade ett jobb åt honom .
jag gav Tom skjuts .
jag fick ett jobberbjudande .
jag blev alldeles upprymd .
jag blev alldeles till mig .
jag fick ett annat jobb .
jag har skaffat ett annat jobb .
jag fick riktigt mycket att göra .
jag blev genomblöt .
jag köpte något gott till dig .
jag fick ditt brev .
jag hade en besvärlig tid .
jag hade det besvärligt .
jag hade det trevligt .
jag kände Tom knappt .
jag känner dig knappt .
jag hatar att komma för sent .
jag avskyr att komma för sent .
jag hatar min bror .
jag avskyr min bror .
jag har ryggont .
jag har ont i ryggen .
jag har ett kontrakt .
jag har en deadline .
jag har huvudvärk .
jag har ont i huvudet .
jag har mycket mera .
jag har en fånge .
jag har en fråga .
jag har en segelbåt .
jag har en gammal bil .
jag har den hemma .
jag har många böcker .
jag har mina skäl .
jag har ingen kommentar .
jag har inga vapen .
jag har några idéer .
jag har lite pengar .
jag har tre barn .
jag måste köpa en .
jag måste hämta Tom .
jag måste få träffa Tom .
jag måste träffa Tom .
jag måste träffa dig .
jag måste sträcka på mig .
jag måste ta det .
jag har arbete att göra .
jag höll Tom i handen .
jag hjälpte Tom en gång .
det tvivlar jag starkt på .
jag hoppas att det hjälper .
jag hoppas att den här fungerar .
jag hoppas kunna lyckas .
jag vet bara inte .
jag hittade dem alldeles nyss .
jag blev just biten .
jag har nyligen flyttat hit .
jag märkte det precis nu .
jag märkte det alldeles nyss .
jag dödade mössen .
det vet jag om .
jag vet om det .
jag känner till hemligheten .
jag vet vem som gjorde det .
jag tycker bättre om Tom .
jag gillar att vara upptagen .
jag gillar utmaningar .
jag tycker om folksånger .
jag gillar den där tröjan .
jag gillar den där skjortan .
jag gillar färgerna .
jag tycker om det här stället .
jag gillar det här stället .
jag tycker om den här platsen .
jag gillar den här platsen .
jag tycker om att vara här .
jag gillar att vara här .
jag gillar din scarf .
jag gillar din halsduk .
jag gillar din sjal .
jag gillar din sjalett .
jag tycker om din scarf .
jag tycker om din halsduk .
jag tycker om din sjal .
jag tycker om din sjalett .
jag tyckte om den där boken .
jag tyckte om den här boken .
jag tappade ett örhänge .
jag förlorade allt .
jag älskar Kalifornien .
jag älskar den där klänningen .
jag älskar den filmen .
jag älskar den scarfen .
jag älskar den halsduken .
jag älskar den sjalen .
jag älskar den sjaletten .
jag älskar den affären .
jag älskar den historian .
jag älskar den sagan .
jag älskar er .
ni har ett jättefint hus .
jag har gjort kaffe åt dig .
jag gjorde kaffe åt dig .
jag har gjort kaffe åt er .
jag gjorde kaffe åt er .
jag kan överleva dig .
jag kan behöva det där .
jag saknar den redan .
jag saknar mina vänner .
jag saknar mitt gamla jobb .
jag saknar dina skämt .
jag har saknat er , barn .
jag måste åka härifrån .
jag behöver Toms hjälp .
jag behöver en dator .
jag behöver en askkopp .
jag behöver en huvudvärkstablett .
jag behöver mer pengar .
jag behöver mina glasögon .
jag behöver lite sömn .
jag behöver lite vatten .
jag behöver de här pengarna .
jag behöver dessa pengar .
jag måste göra det .
jag måste gå vidare .
jag behöver få träffa Tom .
jag behöver träffa Tom .
jag behövde det där jobbet .
jag köper aldrig socker .
jag blir aldrig full .
jag blev aldrig trött .
jag tyckte aldrig om henne .
jag borde gå nu .
jag är skyldig honom 100 yen .
jag spelar fiol .
jag spelade fotboll .
jag läste om det där .
jag tvivlar faktiskt på det .
jag hatar verkligen Tom .
det hoppas jag verkligen inte .
jag tycker verkligen om rött .
jag älskar verkligen Tom .
jag älskar dig verkligen .
jag behöver dig verkligen .
jag kommer ihåg det nu .
jag minns det nu .
jag sa god natt .
god natt , sa jag .
jag sa det fel .
Sväng höger , sa jag .
jag räddade ditt liv .
jag såg Tom tidigare .
jag träffade Tom i kväll .
jag såg Tom i kväll .
jag såg ett flygplan .
jag såg många saker .
jag visste att det där skulle hända .
jag såg meddelandet .
jag visste att det här skulle hända .
jag såg att du tittade .
jag såg dig på utsidan .
jag såg dina fotografier .
jag såg dina foton .
jag skrapade knät .
jag förstår vad problemet är .
jag borde vara där .
jag borde hjälpa Tom .
jag borde tala om det för Tom .
jag sov väldigt bra .
jag sov mycket gott .
jag har ännu tid .
jag har fortfarande tid .
jag pratade för mycket .
jag tror att jag svimmade .
jag tror att jag stannar .
jag tror att det är över .
jag försökte skrika .
jag sa nej till Tom .
jag vände sida .
jag vill ha den här hundvalpen .
jag vill vara här .
jag vill åka tillbaka .
jag vill gå tillbaka .
jag vill träffa Tom .
jag ville ha det bästa .
jag ville ha den bästa .
jag skämdes .
jag hade det trevligt .
jag njöt av det .
han hjälpte till .
jag var på området .
jag var bara rädd .
jag var utmattad .
jag har aldrig varit modig .
jag var på listan .
jag var rätt upptagen .
jag citerade Tom .
jag var verkligen sen .
jag var jättesen .
jag var mycket artig .
jag tittade på tv .
jag var inte alltför upptagen .
jag såg Tom dö .
jag såg på när Tom dog .
jag såg en film .
jag tittade på en film .
jag ska underrätta Tom .
jag ropade efter hjälp .
jag kommer tillbaka snart .
jag är i bilen .
jag kommer att vara ensam .
det gör säkert ont .
jag slår vad om att det gör ont .
jag går och kollar till Tom .
jag ska kolla till Tom .
jag gör det ändå .
jag gör det i alla fall .
jag hämtar mina verktyg .
jag hämtar lite is .
jag hämtar boken .
jag ska hämta boken .
jag går och öppnar .
jag hämtar maten .
jag hämtar gevären .
jag hämtar vinet .
jag går och hämtar dem nu .
jag ordnar en taxi åt oss .
jag går och ser efter .
jag ska gå till skolan .
jag tar någonting att dricka .
jag undersöka det .
jag forska i det .
jag tar jobbet .
jag tar arbetet .
jag ska jobba på det .
jag är också kanadensare .
jag är bra på att köra bil .
jag är frisör .
jag är lite upptagen .
jag är lite öm .
jag är en tålmodig man .
jag är alldeles ensam nu .
jag är helt ensam nu .
jag är ensambarn .
jag är hemskt trött .
jag kommer till dig .
jag är ganska hungrig .
jag är tämligen hungrig .
jag är rätt hungrig .
jag ska skaffa katt .
jag är glad att jag gjorde det .
jag gör det gärna .
jag är glad att vi är överens .
jag kommer att stanna .
jag tänker stanna .
jag är bra på spel .
jag är på dåligt humör .
jag har pyjamasen på mig .
jag är bara en vän .
jag är bara en kompis .
jag chansar bara .
jag är precis som du .
jag är sen till jobbet .
jag är sen till arbetet .
jag är ingen expert .
jag är inte någon expert .
jag ger inte upp .
jag går inte ut .
jag har inte bråttom .
jag är inte välbetald .
det är inte säkert här .
det är inte tryggt här .
jag är inte särskilt upptagen .
jag är gammeldags .
jag har bakjour i dag .
jag är på väg nu .
jag är på g nu .
jag är verkligen ensam .
jag är fruktansvärt upptagen .
jag är din chef nu .
jag har köpt en bil .
jag har en kupong .
jag har en rabattkupong .
jag måste lugna ner mig .
jag måste ta det lugnt .
jag måste plugga .
jag har hört talas om Tom .
är en av er Tom ?
det kunde vara värre .
det är ganska kallt .
den har ingen streckkod .
det måste vara ett tecken .
det låter hälsosamt .
den var inte på rea .
det var inte på rea .
det är en ordbok .
det är en jättebra sång .
det var så länge sedan .
det är hemligt .
det går fint !
det är svårt att säga .
den är i min ficka .
det är i min ficka .
det är bara en dröm .
den är min brors .
det är min brors .
det är ingen hemlighet .
det är inte någon hemlighet .
det är inte färdigt än .
den är inte färdig än .
det är inte klart än .
det är nu eller aldrig .
den ligger på ditt skrivbord .
det ligger på ditt skrivbord .
den ligger på ert skrivbord .
det ligger på ert skrivbord .
den ligger på ditt bord .
det ligger på ditt bord .
den ligger på ert bord .
det ligger på ert bord .
den ligger på din bänk .
det ligger på din bänk .
den ligger på katedern .
det ligger på katedern .
den står på ditt skrivbord .
det står på ditt skrivbord .
den står på ert skrivbord .
det står på ert skrivbord .
den står på ditt bord .
det står på ditt bord .
den står på ert bord .
det står på ert bord .
den står på din bänk .
det står på din bänk .
den står på katedern .
det står på katedern .
den sitter på ditt skrivbord .
det sitter på ditt skrivbord .
det sitter på ert skrivbord .
det sitter på ditt bord .
den sitter på ert bord .
det sitter på ert bord .
den sitter på din bänk .
det sitter på din bänk .
den sitter på katedern .
det sitter på katedern .
det är samma .
det är dags att vi går .
det är dags att vi åker .
det är en våning upp .
håll ett öga på den .
släpp mina armar .
släpp taget om mina armar .
släpp mitt hår .
låt oss göra affärer .
kom så går vi och lägger oss .
låt oss gå och sova .
livet är vackert .
får jag se ditt ID @-@ kort ?
får jag prova den här ?
gå bort från mig .
min hörsel är dålig .
min häst är svart .
mina ben är trötta .
mitt liv är tråkigt .
ingen kan fly .
ingen kan komma undan .
ingen saknas .
ingen litar på Tom .
ingen av oss såg det .
ingen av oss såg den .
nu har jag dåligt samvete .
var nu försiktig .
sitt kvar här nu .
stanna kvar här nu .
vänta lite nu .
vad ska vi göra nu ?
det är klart att han ljög .
Överlappning kan inträffa .
vi ses nästa vecka !
vi ses nästa vecka !
hon kan inte stoppa mig .
hon svor högt .
hon stiger upp tidigt .
hon har en bild .
hon är aggressiv .
hon är inte gift .
hon säljer blommor .
Underteckna på den här raden .
Signera på raden här .
Lukta på den här blomman .
Lös problemet .
någon svarade .
det var någon som svarade .
någon saknas .
någon fattas .
det är någon som saknas .
det är någon som fattas .
prata långsammare .
spindlar spinner nät .
sluta plåga mig .
sluta tjata på mig .
sluta trakassera mig !
sluta trakassera mig .
sluta besvära mig .
säg till Tom att jag är sjuk .
berätta det för Tom .
säg att jag har fel .
berätta för mig om Tom .
säg att det är sant .
berätta din plan för mig .
berätta er plan för mig .
Termiter äter trä .
dörren är låst .
dörrklockan ringde .
maten är färdig .
killen hade en pistol .
hästen är min .
risken är liten .
rummet var mörkt .
världen är ond .
dom talade inte .
de pratade inte .
de talade inte .
de ville ha bevis .
de var perfekta .
de är kannibaler .
de är dyra .
denna bok duger .
den här boken duger .
det här ägget är färskt .
detta är inkorrekt .
det här är inkorrekt .
detta är oriktigt .
det här är oriktigt .
detta är felaktigt .
det här är felaktigt .
den här är jättehäftig .
detta är väldigt lätt .
det här är din hållplats .
det här gör mig arg .
den här är ren .
det här rummet är kallt .
kasta bollen till mig .
Tom åt någonting .
Tom började prata .
Tom började tala .
så kan Tom inte göra .
Tom kan inte göra så .
Tom kan inte göra det .
Tom får inte göra det .
Tom kan inte skada mig .
Tom får inte skada mig .
Tom kan inte se dig .
Tom får inte se dig .
Tom kan inte träffa dig .
Tom får inte träffa dig .
Tom föraktar Mary .
Tom såg det inte .
Tom såg inte det .
Tom dog den dagen .
Tom hade inget val .
Tom är skadad .
Tom har blivit skadad .
Tom hatade sig själv .
Tom hatade spenat .
Tom hatar att dansa .
Tom avskyr att dansa .
Tom hatar att springa .
Tom hatar löpning .
Tom hatar hemligheter .
Tom hatar spindlar .
Tom skadade knät .
Tom är en körgosse .
Tom är sångare i gosskör .
Tom är en flykting .
Tom är en rymling .
Tom är en landsflykting .
Tom är aggressiv .
Tom är alltid varm .
Tom är alltid het .
Tom är vältalig .
Tom är talför .
Tom är förvånad .
Tom är på baren .
Tom är bakom dig .
Tom är trovärdig .
Tom är modig .
Tom är missmodig .
Tom är beslutsam .
Tom är förkrossad .
Tom är diplomatisk .
Tom är missnöjd .
Tom är missbelåten .
Tom håller på att somna .
Tom är illa ute .
Tom är i knipa .
Tom har problem .
Tom är min make .
Tom är min man .
Tom är svarslös .
Tom kommer inte .
Tom är ganska gammal .
Tom är otrogen .
Tom är trolös .
Tom är klarvaken .
Tom är inte sig själv .
Tom sitter inte i fängelse .
Tom är inte i häkte .
Tom sitter inte i häkte .
Tom är inte här uppe .
Tom fortsatte klättra .
Tom gillar det kallt .
Tom tycker om hummer .
Tom gillar att fiska .
Tom tycker om att fiska .
Tom tycker om att sticka .
Tom såg sig omkring .
Tom såg skyldig ut .
Tom ser fantastisk ut .
Tom ser irriterad ut .
Tom ser besvärad ut .
Tom ser ängslig ut .
Tom ser förkrossad ut .
Tom älskade bananer .
Tom fick Mary att gråta .
Tom behöver en tjänst .
Tom kandiderade som borgmästare .
Tom lurade mig .
Tom sjöng för Mary .
Tom visade oss hur .
Tom vill ha hjälp .
Tom vill leka .
Tom vill spela .
Tom var deprimerad .
Tom låg i koma .
Tom kommer att vara här .
Tom kommer nog att tänka om .
Tom förstår nog .
Tom kommer att förstå .
Tom , var är vi ?
prova den där skjortan .
försök att vara i tid .
försök vara i tid .
vänta , skjut inte !
titta på hur jag gör det .
titta hur jag gör det .
kolla hur jag gör det .
vi är de vi är .
vi är inte seriösa .
vi kan båda göra det .
vi kan kolla upp det .
vi kan inte hjälpa dig .
vi kan inte hjälpa er .
vi stänger kl. 19 .
vi stänger 19 .
vi blev stupfulla .
vi hamnade i bråk .
vi satte oss i bilen .
vi hade en bra dag .
vi måste prova det .
vi har inte misslyckats .
vi hoppas på fred .
vi måste betala skatt .
vi satt och väntade .
vi vill ha revansch .
vi vill ha en sak .
vi åkte rakt norrut .
vi åkte till Boston .
vi var väldigt upptagna .
vi var inte roade .
vi ska slutföra den .
vi vann slaget .
vi kommer till det .
vi följer med .
vi är alla släkt .
vi har slut på mjölk .
vi är verkligen upptagna .
vi har nyckeln .
vi måste gömma oss .
vi måste prata .
vilken fantastisk utsikt !
vilken konstig idé !
vad gör vi ?
vad kan Tom göra ?
vad kunde Tom göra ?
vad skulle Tom kunna göra ?
vad visste Tom ?
vad menade Tom ?
vad behövde Tom ?
vad ville Tom ?
vad ville Tom ha ?
vad kände du ?
vad hade du ?
vad menade du ?
vad sjöng du ?
vad gör jag härnäst ?
vad gör jag sen ?
vad ska jag göra sedan ?
vad är jag skyldig dig ?
vad är jag skyldig er ?
vad vet de ?
vad menar de ?
vad gör vi nu ?
vad har Tom sagt ?
vad har Tom sett ?
vad hjälper det ?
vad kallas den ?
vad heter den ?
vad är din idé ?
vad tänker du om det här ?
vad är din uppfattning ?
vad finns i lådan ?
vad är det som luktar ?
vad är det där för lukt ?
vad är det värt ?
vad är det där värt ?
vad är den där värd ?
vad har du hittat ?
var är mina barn ?
var är utgången ?
var ligger utgången ?
var är min chaufför ?
Varifrån kommer den här ?
Varifrån kommer det här ?
Varifrån är den här ?
Varifrån är det här ?
var kommer den här ifrån ?
var kommer det här ifrån ?
var är den här ifrån ?
var är det här ifrån ?
vilken tand gör ont ?
vem kan jag tala med ?
vem kan jag prata med ?
vem gav den till mig ?
vem hjälper dig ?
varför är de här ?
varför ljuger du ?
varför gjorde Tom det ?
varför gjorde hon det ?
varför gör de det ?
varför ge den till mig ?
varför är den inte här ?
varför är det inte här ?
Wow ! vad billigt !
du är i vägen .
du står i vägen för mig .
du är min pappa .
du är min far .
du är en av oss .
du kan parkera här .
du kan lita på honom .
du kan inte rädda mig .
ni kan inte rädda mig .
du kunde ha dött .
du kunde ha stuckit .
ni kunde ha stuckit .
du gjorde ett dåligt jobb .
du gör ett fint jobb .
du gav den till mig .
ni gav den till mig .
ni gav den till oss .
du gav den till oss .
du tappade tilltron till mig .
du ser tveksam ut .
ni ser tveksamma ut .
du ser bekant ut .
du får parkera här .
du måste hjälpa henne .
ni måste hjälpa henne .
du behöver koppla av .
du borde veta .
du är skyldig mig en öl .
ni är skyldiga mig en öl .
du pratar för mycket .
du är aggressiv .
ni är aggressiva .
du kväver mig .
du håller på att kväva mig .
du kan gå .
du sitter på min plats .
du ljuger ju bara .
ni ljuger ju bara .
du har rätt , Tom .
ditt hus är stort .
ert hus är stort .
ett barn är försvunnet .
det är en vakt på utsidan .
det är mycket som har hänt .
allt är lugnt igen .
vi är alla upptagna .
är jag fånig ?
stör jag dig ?
håller vi tidtabellen ?
är du buddist ?
är du buddhist ?
är du en fånge ?
är du svårt skadad ?
Skyller du på mig ?
är ni två fulla ?
är ni båda fulla ?
har du det bra ?
är ni beväpnade ?
känner ni varandra väl ?
är ni galna ?
är ni färdiga ?
är du hungrig ännu ?
är ni hungriga ännu ?
gör du narr av mig ?
är du verkligen Tom ?
är du fortfarande upptagen ?
är ni två hungriga ?
är dina ögon öppna ?
bananer är gula .
öl innehåller humle .
Attans , det var nära .
frukosten är färdig .
ta Tom med dig .
köp lågt , sälj högt .
kan jag låna en penna ?
får jag låna din ?
kan jag räkna med Tom ?
kan jag göra det själv ?
får jag göra det själv ?
kan jag få en kudde ?
kan jag få pengarna tillbaka ?
kan jag få en tatuering ?
kan jag gömma mig här ?
kan jag gömma mig här inne ?
får jag förhöra Tom ?
får jag ställa frågor till Tom ?
kan jag säga det högt ?
får jag sitta med Tom ?
kan jag sitta med Tom ?
får jag tala med Tom ?
får jag prata med Tom ?
kan jag ta en paus ?
kan jag tala om för Tom varför ?
kan man lita på Tom ?
har vi råd med det där ?
har vi råd med det här ?
kan vi sätta igång ?
kan du ordna det ?
kan du förlåta oss ?
kan du hålla tyst ?
kan du förhindra det ?
kan du skydda mig ?
kan du skydda oss ?
kan du bevisa det ?
kan du se någon ?
kan du gå ännu ?
kan du lita på dem ?
kan du inte se det ?
kolla in den här .
barn behöver kärlek .
städa upp den här röran .
kom tillbaks om en dag .
kom tillbaks om ett dygn .
kom hit en sekund .
kom och hälsa på oss snart .
Behärska er .
kan Tom ha fel ?
kan vi gå nu ?
kan vi beställa nu ?
ta itu med det senare .
sa jag för mycket ?
trodde Tom på det ?
har Tom ätit middag ?
åt Tom middag ?
jobbade Tom där ?
var det någon som saknade mig ?
fick du fast dem ?
tyckte du om det där ?
njöt du av det där ?
kidnappade du Tom ?
var det du som kidnappade Tom ?
var det du som mördade Tom ?
har du underrättat Tom ?
har du meddelat Tom ?
målade du det här ?
sov du här ?
gjorde du anteckningar ?
hörde du mig inte ?
hörde ni mig inte ?
middagen var toppen .
ser jag ut som Tom ?
behöver jag en orsak ?
måste jag skynda mig ?
är jag skyldig dig pengar ?
är det kakor jag känner doften av ?
gör som jag säger åt dig .
säljer de böcker ?
misstänker de mig ?
tar ni emot dricks ?
hör du hemma här ?
känner du dig hungrig ?
har du en kopia ?
har du någon legitimation ?
har du tillräckligt ?
gillar du Mozart ?
tycker du om Mozart ?
gillar du ost ?
tycker du om städer ?
tycker du om storstäder ?
tycker du om kaffe ?
tycker du om att vandra ?
tycker du om att gå på vandring ?
tycker du om robotar ?
tycker du om lax ?
tycker du om skolan ?
gillar du skolan ?
tycker du om sommaren ?
tycker du om sommar ?
saknar du Boston ?
behöver du hjälp ?
behöver du den nu ?
behöver ni den nu ?
spelar du squash ?
spelar du tennis ?
kommer du ihåg oss ?
känner du att det luktar rök ?
dansar du fortfarande ?
vill du ha lift ?
vill du ha skjuts ?
läkare räddar liv .
behöver Tom hjälp ?
stör det dig ?
Involverar det mig ?
Behagar det dig ?
gör det fortfarande ont ?
fungerar den ännu ?
jobbar hon hårt ?
betyder det ja ?
var inte arg på mig .
bli inte paranoid .
bli inte överkörd .
bli inte så arg .
ge inte bort den .
Skänk inte bort den .
avslöja det inte .
släpp mig inte .
släpp inte taget om mig .
gör honom inte besviken .
Ställ inte till en scen .
prata inte strunt .
tacka mig inte än .
ner med kungen !
drick med mig , Tom .
till och med Tom tycker det .
alla fick panik .
alla satt sig ned .
alla satt sig ner .
alla tvekade .
alla väntar .
alla står och väntar .
allt förändrades .
allt förändras .
allt slutade .
allt är fel .
ursäkta mig ett ögonblick .
ursäkta mig en sekund .
förklara det för mig .
fyll i det här formuläret .
ge eld på mitt kommando .
glöm att jag sa det där .
glöm vad jag sa .
hämta lite vatten åt Tom .
kolla in den här .
hämta en shot av det här .
gå bort från det där .
gå till era platser .
hämta lite kaffe åt mig .
kom ner från mitt tak .
kom hit , Tom .
gör er redo för avfärd .
gör dig redo för avfärd .
gör dig av med pistolen .
hämta din rock , Tom .
skaffa en egen lägenhet .
ge Tom allting .
ge Tom lite utrymme .
ge din sittplats till Tom .
ge mig ett exempel .
ge mig min andel .
ge mig lite pengar .
ge mig lite plats .
ge mig lite vatten .
ge mig den där .
ge mig rapporten .
ge mig dina händer .
ge mig din kniv .
ge mig din tröja .
gör det nu bara .
gå och ta en titt .
gå och tala med Tom .
gå runt den vägen .
gå och fråga din far .
gå och lägg dig igen nu .
gå och borsta håret .
gå och hämta lite handdukar .
gå hem och byt kläder .
gå upp för den här trappan .
gå och vänta i bilen .
gissa vad jag hittade .
slå in spiken .
ge mig den där kvasten .
ge mig brevet .
ge mig tången .
vänta en sekund .
stanna kvar en sekund .
hårt arbete lönar sig .
har Tom fått sparken ?
har jag missat mycket ?
ha en bra sommar .
se dig runt .
ta ett glas till .
ha så kul i Boston .
ha så roligt i Boston .
har du varit fattig ?
har du glömt ?
har du ätit lunch ?
har du läst det här ?
har du sett det här ?
han kom fram i tid .
har tråkar ut allihopa .
han dog i sin säng .
han lyssnar inte .
han känner inte mig .
han klarade det till slut .
han glömde hennes namn .
han glömde det igen .
han kom förbi mig .
han var tvungen att gå dit .
han har en vit hund .
han höll andan .
han är en dålig chaufför .
han är alltid glad .
han har alltid rätt .
han är inte läkare .
han spelar golf .
han är segraren .
han behöll hatten på .
han låg på rygg .
han lever i lyx .
han älskar att resa .
han kan vara ett geni .
han föste iväg henne .
han skapade ett prejudikat .
han rakade huvudet .
han väntade på sin tur .
han var riktigt kall .
han tog en promenad .
han är en drama queen .
han är redan en man .
han är duktig med kort .
han är inte ett olydligt barn .
hjälp ! jag drunknar !
här kommer Tom nu .
här är ett exempel .
här är lite vatten .
här har du lite vatten .
här , ta en drink .
här , ta någonting att dricka .
här , smaka en bit .
Hallå , öppna dörren .
Hallå där , lägg tillbaka den där .
hans fötter är smutsiga .
vänta en sekund .
skulle det smaka med lite te ?
vad tycker du om den här ?
hur noggrann är den ?
hur pass noggrann är den ?
hur mår de andra ?
hur stor kommer den att vara ?
hur kan jag hjälpa Tom ?
hur kan jag stoppa Tom ?
hur kan vi göra det ?
hur kan du laga den ?
hur bra kände ni varandra ?
hur skulle jag kunna glömma ?
hur kunde Tom veta det ?
hur betedde Tom sig ?
hur kom Tom in ?
hur tog sig Tom in ?
hur tog Tom sig in ?
hur har Tom fått den ?
hur gick det , Tom ?
hur åkte de ?
hur gjorde vi det ?
hur missade vi det ?
hur flydde du ?
hur lyckades du fly ?
hur ska jag tacka dig ?
hur ska vi hitta Tom ?
hur hittar vi Tom ?
hur hittar vi ut ?
hur ska vi stoppa Tom ?
hur känns det ?
hur känns det där ?
hur ser det här ut ?
hur långt kan du gå ?
hur långt gick du ?
hur svårt kan det vara ?
hur känner Tom sig ?
hur mår din far ?
hur stora är de ?
hur länge sedan är det ?
vad kostar en öl ?
hur gammal är Tom nu ?
hur säkert är Brasilien ?
hur var det igår kväll ?
hur var baletten ?
hur var flygresan ?
hur var din kväll ?
hur skulle Tom veta det ?
hur skulle du veta ?
hur kom du hit ?
hur känner du dig ?
hur mår din patient ?
jag håller fullständigt med .
jag beundrar Tom mycket .
jag ljuger nästan aldrig .
jag har redan sagt det till dig .
jag är enda barnet .
jag är inte för trött .
jag kom för sent .
jag frågade vem han var .
jag åt alldeles för mycket .
jag tror på allt det där .
jag tog med mig Tom hit .
jag förde Tom hem .
jag brände pappret .
jag brände papperet .
jag brände soporna .
jag kan ordna det .
jag kan vara artig .
jag kan övertalas .
det kan jag tro på .
jag kan ta itu med det .
jag kan köra själv .
jag kan förklara det där .
det kan jag förklara .
jag kan förklara det här .
jag kan knappt stå .
jag kan hjälpa dig .
jag kan föreställa mig det .
jag kan leva med det .
jag kan stå ut med det .
jag kan betala tillbaka .
det kan jag respektera .
jag inser det nu .
jag kan tala med Tom .
jag kan inte tillåta det .
jag kan inte bryta mig loss .
jag kan inte bryta mig fri .
jag kan inte bara gå .
jag tål inte golf .
jag kan inte förstå .
jag samåker med Tom .
jag bytte skjorta .
jag dubbelkollade det .
jag kollade det två gånger .
jag kontrollerade det två gånger .
jag kollade datumet .
jag kollade med Tom .
jag skulle kunna ha rätt .
det kan vara till hjälp .
det skulle sitta fint med en öl .
jag kunde behöva lite hjälp .
jag kunde ha drunknat .
jag kunde ha sagt nej .
jag knäckte koden .
jag kräver sanningen .
jag gjorde det helt själv .
jag gjorde det frivilligt .
jag gjorde mitt arbete väl .
jag överraskade verkligen Tom .
det visste jag inte .
jag rörde inte Tom .
jag ville inte ha mjölk .
jag har inget jobb .
jag har ingen vodka .
jag förstår inte .
jag drack kaffet .
jag tyckte om att simma .
jag förväntar mig din hjälp .
jag känner en smärta här .
jag känner mig så hjälplös .
jag känner mig väldigt skyldig .
jag känner mig väldigt stark .
jag föll av min cykel .
jag kände mig skyldig .
jag kände mig väldigt sömnig .
jag kände mig väldigt illa till mods .
jag antog det .
jag vann över Tom till slut .
jag tvingade honom att gå .
jag glömde min plånbok .
jag hittade lite pengar .
jag hittade din dagbok .
jag fann din dagbok .
jag gav Tom mitt ord .
jag gav upp för tidigt .
jag lovar .
jag missförstod allting .
jag har gjort mig fin i håret .
jag fick ditt meddelande .
jag fick en uppenbarelse .
det har varit en hemsk dag .
jag har haft en hemsk dag .
jag hade lite problem .
jag fick den där känslan .
jag simmar nästan aldrig .
jag hatar min dator .
jag hatar min rumskompis .
jag hatar de här orden .
jag har några idéer .
jag har ett bra arbetslag .
jag har en bra besättning .
jag har ett jättebra jobb .
jag har ett jobb att göra .
jag har en lista här .
jag har hittat ett jobb .
jag har en begäran .
jag har en med mig .
jag har fakturan .
jag har biljetterna .
jag måste åka hem .
jag måste ta mig hem .
jag måste veta det nu .
jag måste repetera .
jag måste säga det här .
jag måste sätta mig .
jag måste sätta mig ner .
jag måste ge mig i väg .
jag har två biljetter .
jag har vad jag behöver .
jag har vad jag vill ha .
jag hörde Tom skrika .
jag gömde den någonstans .
jag hoppas att det är sant .
jag hoppas att det stämmer .
jag hoppas kunna vara med .
jag hoppas att vi slår Tom .
jag hoppas att vi kan hjälpa .
jag hoppas att vi hittar Tom .
jag hoppas att vi finner Tom .
jag hoppas att du tycker om mig .
jag skadade min vänstra arm .
jag har för avsikt att använda den .
jag bjöd hem Tom .
jag lånade den precis .
jag lånade den bara .
jag lånade den just .
jag köpte den här nyss .
jag kan bara inte sova .
jag kan inte sova bara .
jag känner mig bara dum .
jag har nyligen förlovat mig .
jag ville bara ha pengar .
jag behöll tröjan .
jag kände din far .
jag kände din fader .
jag kände din pappa .
jag känner bra till Boston .
jag vet att Tom fuskade .
jag kan min sak .
jag vet vad jag vill .
jag vet vad jag vill ha .
jag vet att du är upptagen .
jag vet att ni är upptagna .
jag känner din mamma .
jag känner din mor .
jag tycker om koreansk mat .
jag gillar Tom redan .
jag gillar fjärilar .
jag tycker om fjärilar .
jag gillar serieböcker .
jag tycker om kapplöpningar .
jag tycker om hallon .
jag gillar den personen .
jag gillar den här gitarren .
jag gillar att vara ensam .
jag tycker om tv @-@ spel .
jag gillade den där filmen .
jag gillade den filmen .
jag gillade din historia .
jag tyckte om din historia .
jag tappade bort mitt häfte .
jag älskar utmaningar .
jag älskar äppeljuice .
jag älskar män med skägg .
jag älskar den där tatueringen .
den där tatueringen är superfin .
jag älskar de där skorna .
jag gjorde den här själv .
jag klarar mig bara fint .
jag träffade honom nyligen .
jag saknar Tom redan .
jag saknar Tom så mycket .
jag behöver en sekreterare .
jag behöver ett kuvert .
jag behöver en timme ledigt .
jag behöver en till .
jag behöver säkra bevis .
jag behöver deras namn .
jag måste motionera .
jag måste mata Tom .
jag måste få veta .
jag måste åka dit .
jag måste hjälpa Tom .
jag måste få veta varför .
jag måste berätta det för Tom .
jag behöver ditt nummer .
jag tvivlade aldrig på det .
jag åkte aldrig fast .
jag gjorde aldrig Tom illa .
jag rörde den aldrig .
jag bär aldrig kostymer .
jag spelar tv @-@ spel .
jag föredrar låga klackar .
jag släckte elden .
jag läste din rapport .
jag hatar verkligen det här .
jag tyckte verkligen om dig .
jag saknar dem verkligen .
jag behöver verkligen det här .
det här behöver jag verkligen .
jag borde faktiskt gå .
jag vill verkligen ha den här .
jag vill verkligen ha det här .
jag träffade nyligen Tom .
jag gick i pension vid sextio .
jag springer två gånger i veckan .
jag sparar mina kvitton .
jag såg bilderna .
jag såg dem kyssas .
jag såg vad Tom gjorde .
jag såg vad du gjorde .
jag borde göra mig färdig .
jag borde gå och byta om .
jag borde veta det .
jag borde stanna här .
jag borde ta den här .
jag borde ha stannat .
jag skulle ha stannat .
jag log för mig själv .
jag vill fortfarande gå .
jag vill fortfarande åka .
jag vill fortfarande fara .
jag föreslår att du duckar .
jag föreslår att du gömmer dig .
jag tror att jag gillar dig .
jag tycker att det är galet .
jag tror att det hjälper .
jag tror att vi är vilse .
jag tror att vi står på tur .
jag tror vi står på tur .
jag tänkte på det .
jag trodde att du slutade .
jag trodde att du slutat .
jag följde ditt råd .
det kan jag helt och hållet förstå .
jag vill ha en advokat .
jag vill träffa Tom .
jag ville byta om .
jag ville förändras .
jag var ironisk .
jag var hövlig .
jag kände mig deppig .
jag läste bara .
jag retades bara .
jag retades bara lite .
jag skämtade bara .
jag retades bara .
jag var stolt över Tom .
jag var ganska hungrig .
jag sov djupt .
jag blev tillsagd att hjälpa .
jag var väldigt självisk .
jag jobbade sent .
jag var inte ens här .
jag tittar på tv .
jag gick till banken .
jag ska skydda dig .
jag önskar att jag hade vetat .
jag arbetade på en bondgård .
det skulle jag tycka om .
jag kunde vara med på det .
jag kunde ställa upp på det .
jag borde nog också gå .
jag är vid mitt skrivbord .
du hittar mig vid mitt skrivbord .
jag ska köpa en ny .
jag bjuder dig på lunch .
jag ska göra som du säger .
jag ska äta äpplet .
jag hämtar den själv .
jag hämtar det själv .
jag ska göra mig färdig nu .
jag ska göra mig av med den .
jag hämtar notan .
jag ska hämta en pistol åt dig .
jag hämtar din rock .
jag hämtar din kappa .
jag hämtar din jacka .
jag går ut på en promenad .
jag går och hämtar den nu .
jag går och hämtar det nu .
jag går och hämtar min bil .
jag åker i natt .
jag åker i kväll .
jag far i natt .
jag far i kväll .
jag kommer att sakna er alla .
jag skall läsa boken .
jag ska läsa boken .
jag dukar .
jag kan gå i god för Tom .
jag är lite galen .
jag är lite tidig .
jag är lite skakig .
jag är fotograf .
jag ska strax gå .
jag är rädd för hundar .
jag är också lärare .
jag är en gammal man nu .
jag är lika lång som du .
jag är lealös .
jag känner mig hungrig .
jag börjar bli hungrig .
jag är glad att jag har träffat dig .
jag är glad att Tom är okej .
jag är glad att det fungerade .
jag är glad att vi pratades vid .
jag är glad att vi väntade .
jag ska ta en joggingrunda .
jag klarar mig .
jag ska göra det .
jag ska studera .
jag följer med Tom .
jag är bra på mitt jobb .
jag gör det gärna .
jag gör det gladeligen .
jag är här ensam .
jag håller på att bli galen .
jag är inte död , eller hur ?
jag är ju inte död , eller hur ?
jag är inte bra på det .
jag är inte lycklig här .
jag är inte intresserad .
jag är inte arg på dig .
jag sticker till gymmet .
jag är verkligen försiktig .
jag är verkligen noggrann .
jag är led på skolan .
jag är less på skolan .
jag är utled på skolan .
jag är så generad .
jag är dubbelt så gammal som du .
jag är lite låg .
jag är deppig .
jag har pengarna .
jag måste bege mig nu .
jag har blivit bättre .
jag tycker också om godis .
är Tom kristen ?
är det någon här inne ?
är det tillräckligt ?
är den här platsen upptagen ?
är inte Tom med dig ?
är inte Tom med er ?
den måste vara där .
det är måndag i dag .
det slutade bra .
det var mitt nöje .
det var bara ett skämt .
det var inte på ovanvåningen .
det får vänta .
det måste vänta .
det är ett stort företag .
det är ett villospår .
det är en avledningsmanöver .
det kommer att regna .
det måste vara nu .
den står i garaget .
den är i garaget .
det är bara en teori .
det är inget misstag .
det är inget problem .
det är inte något problem .
det är inte viktigt !
det är inte mitt val .
det är inte så lite .
det är inte så djupt .
den är inte där nu .
det är inte där nu .
det är inte upp till dig .
det är inte upp till er .
det regnar fortfarande .
det är den andra .
det är fel .
gör bara som jag gjorde .
gör bara som jag säger .
gör ett försök bara .
ge den till mig bara .
sitt och slappna av bara .
sitt och koppla av bara .
sätt dig ned bara , Tom .
sätt dig ner bara , Tom .
Släng iväg den bara .
kasta den bara .
håll dig ur min väg .
håll er ur min väg .
kunskap är makt .
låt mig prata med Tom .
låt mig tala med Tom .
vi ger det ett försök .
kom så äter vi lunch .
kom så går vi hem , Tom .
kom så åker vi hem , Tom .
vi går hem , Tom .
vi åker hem , Tom .
låt oss anordna en fest .
vi släpper det bara .
vi släpper den bara .
kan vi inte bara säga ja ?
vi säger bara ja .
vi fortsätter leta .
vi fortsätter titta .
du , jag måste gå .
Mary är attraktiv .
får jag titta på tv nu ?
gå lite bakåt .
mina väskor är packade .
min familj är liten .
mina händer var fulla .
mitt hjärta är brustet .
min brevlåda är full .
min näsa är för stor .
min plan fungerar .
mitt rum vetter mot öst .
ge aldrig upp hoppet .
ingen är odödlig .
ingen är oskyldig .
ingen får avlägsna sig .
ingen såg någonting .
ingen hjälpte till .
ingen var med mig .
ingen köper det .
ingen köper den .
ingen behöver veta .
det är ingen som bor där .
inget saknas .
nu vill jag vila .
nu har du din chans .
Ligg nu bara stilla .
Ligg nu bara still .
vänta en minut nu .
okej , jag fattar .
ur vägen , pojk .
be för oss allihopa .
råttor förökar sig fort .
kom genast tillbaka .
Återvänd genast .
Återvänd till skeppet .
spara det till senare .
hon kan inte stoppa mig .
hon har solglasögon .
hon hörde honom sjunga .
hon åkte till Paris .
han bor i Kyoto .
hon bor i Kyoto .
hon plockade blommor .
hon vill dansa .
borde vi berätta för Tom ?
så vad gjorde du ?
vatten , tack .
lite vatten , tack .
håll dig borta från Tom .
stanna här med Tom .
stanna , annars skjuter jag .
sluta prata med mig .
sluta upp med det där tramset .
ta ut soporna .
ta bort lådan .
hälsa till Tom .
hälsa Tom att jag är färdig .
säg till Tom att jag är färdig .
säg till Tom att jag är ledsen .
säg hej till Tom från mig .
säg vad vi ska göra .
den där dockan är skrämmande .
det var svårt .
det var poängen .
det var din idé .
det vore oförskämt .
det skulle vara oförskämt .
det får duga .
det är allt du får .
det är allt ni får .
det där är allt du får .
det där är allt ni får .
det där är en av mina .
den där är en av mina .
det är oviktigt .
det är där jag sitter .
äpplena är stora .
pojken hoppar .
klockan är två .
jag bjuder på kaffet .
Kråkan flög iväg .
hunden hoppar .
dörren är låst .
Dörrhandtaget gick sönder .
tjejen är ensam .
flickan är ensam .
isen smälter .
köttet är djupfryst .
Mjölken surnade .
kjolen är grön .
spindeln är död .
sommaren är över .
telefonen ringde .
vattnet är rent .
fönstret är öppet .
det finns en buss här .
det är en buss här .
det är en gasläcka .
det här är mina byxor .
de ser alla glada ut .
de kan inte stoppa oss .
de äter choklad .
de fick en stor en .
de ser förvirrade ut .
de ser bekanta ut .
de ser så lyckliga ut .
de ser så glada ut .
de verkar så lyckliga .
de verkar så glada .
de blev mördade .
de mördades .
de simmade .
de har haft ett snack .
den här boken är tung .
den här pojken är min son .
den här stolen är ful .
den här kostar ingenting .
det här är en dålig idé .
det här är en dålig plan .
det här är till stor hjälp .
det här är en busshållplats .
det här är ett bra jobb .
det här är allt jag har .
det här är allt jag behöver .
det här är allt jag vill ha .
det här är omöjligt .
detta är omöjligt .
detta är skandalöst !
det här är riktigt illa .
det här är löjligt !
det här är väldigt billigt .
den här är väldigt billig .
det här är väldigt färskt .
det här är inte rätt .
det här är inte korrekt .
det här är inte riktigt .
de här pengarna är mina .
den här är större .
den här är från mig .
den här är inte bra .
det här borde hjälpa .
den här soppan är jättegod .
det där är mina skor .
vi har tiden på vår sida .
Tom svimmade nästan .
Tom åt upp ditt godis .
Tom blev ängslig .
Tom spelar på hästar .
Tom sjukanmälde sig .
Tom hör dig inte .
Tom kan inte höra dig .
Tom kan inte skada dig .
Tom kan inte ställa sig upp .
Tom kan inte stå upp .
Tom skulle kunna vara en polis .
Tom gav inte upp .
Tom berättade inte det för mig .
Tom hittade bevis .
Tom satte sig i bilen .
Tom blev väldigt arg .
Tom hängde sig .
Tom har svimmat .
Tom har tuppat av .
Tom har kolat av .
Tom har kort hår .
Tom måste gå hem .
Tom hatar barn .
Tom avbröt mig .
Tom är en bra grabb .
Tom är en mäktig man .
Tom är en smart grabb .
Tom är sociopat .
Tom ska precis gå .
Tom är äventyrlig .
Tom är vid dörren .
Tom är karismatisk .
Tom kommer tillbaka .
Tom är tävlingsinriktad .
Tom är tävlingslysten .
Tom är omtänksam .
Tom är samarbetsvillig .
Tom är missnöjd .
Tom är olydig .
Tom är nedstämd .
Tom är mållös .
Tom är häpen .
Tom är förbluffad .
Tom är förstummad .
Tom är enastående .
Tom är erfaren .
Tom har aldrig fel .
Tom är på lastkajen .
Tom är på lastningsplatsen .
Tom är väldigt snabbt .
Tom är jättesnabb .
Tom är där .
Tom är fortfarande vid liv .
Tom är omöjlig att hindra .
Tom är omöjlig att stoppa .
Tom är ohejdbar .
Tom är din vän .
Tom är inte något hot .
Tom är inte därinne .
Tom är inte som du .
Tom är inte likadan som du .
Tom är inte min fiende .
Tom dök precis upp .
Tom dök bara upp .
Tom var medveten om riskerna .
Tom skrattade högt .
Tom tycker om simning .
Tom haltar lätt .
Tom såg irriterad ut .
Tom tittade på Mary .
Tom såg förbryllad ut .
Tom såg villrådig ut .
Tom såg häpen ut .
Tom såg frågande ut .
Tom ser orolig ut .
Tom ser upphetsad ut .
Tom ser upprörd ut .
Tom ser förskräckt ut .
Tom såg förbryllad ut .
Tom ser förvirrad ut .
Tom ser konfys ut .
Tom ser konfunderad ut .
Tom ser omtumlad ut .
Tom ser ångerfull ut .
Tom ser bekant ut .
Tom ser ut som du .
Tom ser lättad ut .
Tom ser så lycklig ut .
Tom ser så glad ut .
Tom fick Mary att sluta .
Tom har kanske rätt .
Tom måste hjälpas .
Tom fick slut på bensin .
Tom satt bredvid mig .
Tom säger att han är upptagen .
Tom verkar stressad .
Tom skickade mig ett meddelande .
Tom skakade på huvudet .
Tom borde vara här .
Tom tog någonting .
Tom ville hämnas .
Tom vill ha bevis .
Tom vill ha vår hjälp .
Tom vill ha dig tillbaka .
Tom var otrolig .
Tom var ofattbar .
Tom var fantastisk .
Tom var väldigt modig .
Tom kommer inte att vara redo .
Tom kommer inte att vara färdig .
Tom kommer inte att skada dig .
Tom skrek åt Mary .
Tom skrek på Mary .
Toms hund ställde sig upp .
Toms näsa var röd .
Tom är inte färdig .
Tom är inte klar .
Tom är inte hemma än .
försök att inte bli sen .
stäng av vattnet .
blev någon dödad ?
att titta på tv är roligt .
det är roligt att titta på tv .
det är kul att titta på tv .
vi grät mycket allihopa .
alla måste vi dö .
vi är vad vi är .
vi kom för att träffa dig .
vi kan alla göra det här .
vi kan lita på Tom .
vi fattar vinken .
vi kan inte dödas .
vi får inte dödas .
vi kan inte göra det nu .
vi får inte göra det nu .
vi gör som vi vill .
vi odlar vete här .
vi hade ett stort gräl .
vi hade ett stort bråk .
vi hade det trevligt .
vi hade det trevligt .
vi hade en tuff dag .
vi har haft en tuff dag .
vi fick hjälpa Tom .
vi har inga hemligheter .
vi måste göra det där .
vi måste göra det här .
du måste springa nu .
vi lyssnar på musik .
vi behöver Toms hjälp .
vi behöver en ny plan .
vi måste vara säkra .
vi måste hitta den .
vi måste hitta det .
vi måste testa den .
vi spelade baseboll .
vi borde ringa Tom .
vi tog en promenad .
vi var alla rädda .
vi var väldigt lyckliga .
vi var väldigt glada .
vi var unga då .
vi klarar oss .
vi kommer att klara oss .
vi skaffar nya .
vi får nya .
vi ger tillbaka den .
vi ger tillbaka det .
vi giver tillbaka den .
vi giver tillbaka det .
vi ska ha fest .
vi måste vänta .
vi kommer att behöva vänta .
vi kommer att måsta vänta .
vi får det att fungera .
vi har pratat färdigt .
vi kommer att försöka .
vi är goda vänner .
vi finns här för dig .
vi är utom fara .
vi är inte ett par .
vi är inte döda än .
vi är sena .
vi är klara här .
vi är väldigt nöjda .
vi är väldigt belåtna .
vi har kommit för att hjälpa till .
vi har en kvar .
vi måste skynda oss .
vi måste åka härifrån .
var de bra ?
var de med dig ?
stod ni två nära varandra ?
vilken rörig dag .
vilken smart idé !
vad är jag här för ?
vilken förfärlig röra !
vilken ful klänning !
vad blev det av Tom ?
vad kan vi förvänta oss ?
vad har du att erbjuda ?
vilket ackord är det ?
vad kan det betyda ?
vad kunde det vara ?
vad kunde det här vara ?
vad beställde Tom ?
vad svarade Tom ?
vad tyckte Tom ?
vad ansåg Tom ?
vad skrev Tom ?
vad svarade hon ?
vad betydde det ?
vad betydde det där ?
vad tog de ?
vad ville de ?
vad tog du med dig ?
vad hade du med dig ?
vad lärde du dig ?
vad beställde du ?
vad spillde du ?
vad stal du ?
vad var det du stal ?
vad tyckte du ?
vad tittade du på ?
vad ska jag kalla dig ?
vad säger jag till Tom ?
vad ska jag säga till Tom ?
vad tycker de ?
vad anser de ?
vad är vi skyldiga Tom ?
hur mycket tar du ?
vad har hon ?
vad annat finns det ?
vilken våning är jag på ?
vad hände sen ?
vad hände sen ?
vad hände sedan ?
och om han har fel ?
vad är mitt saldo ?
vad är det där borta ?
vad är det som luktar ?
vad är det där för lukt ?
vad är det där för ljud ?
vad är det som låter ?
vad är det där för någonting ?
vad är det här för någonting ?
vilken station är det här ?
vilken station är detta ?
vad skulle ha veta ?
varför dröjer Tom ?
vad uppehåller Tom ?
vad är avbrottet ?
vad är problemet ?
vad är det med Tom ?
när kan jag flytta in ?
när kan jag träffa Tom ?
när vill vi ha det ?
när vill vi ha den ?
när använder du den ?
när börjar det ?
när kommer Tom ?
när börjar det ?
när är begravningen ?
var är mina stövlar ?
var är nycklarna ?
var är barnen ?
var är du , Tom ?
var satte jag den ?
var bodde du någonstans ?
var bodde du ?
var bodde ni ?
var ska jag stiga av ?
var ska jag anmäla mig ?
var ligger hotellet ?
var är ditt rum ?
vart ska vi gå ?
var är Tom född ?
vart är smöret ?
vem gav den till dig ?
vem är din advokat ?
vem är er advokat ?
vem vill ha den här ?
vem vill ha det här ?
vem vill slåss ?
vem är det som överdriver ?
vem är med Tom nu ?
vem är din lärare ?
vems rum är det här ?
varför kan inte Tom tala ?
varför kan inte Tom prata ?
varför kan du inte komma ?
varför frågade du mig ?
varför behöver jag hjälp ?
varför gör du sådär ?
varför gör du såhär ?
varför tycker du om det ?
varför vill du ha den ?
varför vill du ha det ?
varför slutar du inte ?
varför slutar ni inte ?
varför är Tom så upptagen ?
varför är han så tyst ?
varför är inte Tom här ?
varför var du där ?
du sitter på min plats .
du är på min plats .
du kan också göra det .
du kan inte backa ur .
du får inte backa ur .
du kan inte hoppa av .
du får inte hoppa av .
du får inte smita .
du kan inte skylla på mig .
du får inte skylla på mig .
du får inte ringa Tom .
du får inte skada Tom .
du kan inte skada Tom .
ni får inte skada Tom .
ni kan inte skada Tom .
du kan inte lämna mig .
du får inte lämna mig .
ni får inte lämna mig .
du kan inte sluta nu .
du får inte sluta nu .
ni får inte sluta nu .
ni kan inte sluta nu .
det sade du inte .
du skrämmer mig inte .
ni har rätt .
ditt hår ser hemskt ut .
du måste stiga upp .
du måste gå nu .
du måste se det .
du har två bollar .
du kan reglerna .
du kanske har rätt .
du har kanske rätt .
du får inte röka .
ni får inte röka .
du behöver ny bil .
du behöver en ny bil .
du behöver en ny .
du måste gå nu .
du verkar förvånad .
du var dålig på det .
du låg i koma .
du kommer inte att tycka om Tom .
du kommer inte att gilla Tom .
ni kommer inte att tycka om Tom .
ni kommer inte att gilla Tom .
ni är alla bjudna .
du är karismatisk .
ni är karismatiska .
du är tidig igen .
ni är tidiga igen .
du är gift nu .
ni är gifta nu .
du hjälper inte till .
ni hjälper inte till .
du är så paranoid .
ni är så paranoida .
du är fortfarande ung .
du har en timme på dig .
du har en timma på dig .
ni har en timme på er .
ni har en timma på er .
din andedräkt stinker .
hos dig eller hos mig ?
&quot; lita på mig &quot; , sade han .
en tupplur vore bra .
allt jag kan göra är försöka .
låt mig förklara .
ska jag bli utbytt ?
stör jag dig ?
stör jag er ?
gör jag det rätt ?
Inbillar jag mig det här ?
svara mig genast .
vill någon ha en öl ?
det kan vem som helst se .
är de alla starka ?
är de fortfarande här ?
är det där nya skor ?
är det där dina väskor ?
är vi nästan framme ?
är du polis ?
är du polisman ?
är du nästan klar ?
kommer du tillbaka ?
kommer du , Tom ?
är du från Boston ?
tänker du följa med ?
gråter ni ?
försöker du blåsa mig ?
är ni hungriga , barn ?
ljuger du för mig ?
finns du på Facebook ?
har du Facebook ?
är du på semester ?
är ni från vettet ?
är du verkligen upptagen ?
är du verkligen klar ?
är du helt säker ?
är du fortfarande ensam ?
är du fortfarande yr ?
är du så dum ?
är ni två släkt ?
tittar du på mig ?
frukosten är serverad .
ta med dig din verktygsback .
får jag bjuda dig på lunch ?
kan jag ringa upp dig ?
kan jag komma med Tom ?
kan jag komma med dig ?
kan jag göra det för dig ?
kan jag göra det åt dig ?
får jag ta en bild ?
kan jag få ett kvitto ?
får jag ge den här till dig ?
kan jag gå och lägga mig nu ?
kan jag också få en ?
kan jag få listan ?
kan jag åka med dig ?
kan jag säga en sak ?
kan jag träffa dig senare ?
kan jag stanna och hjälpa till ?
kan jag ta med mig Tom hem ?
får jag följa dig hem ?
kan någon hjälpa mig ?
kan någon höra oss ?
kan vi göra någonting ?
kan vi bara gå hem ?
kan vi prata franska ?
kan vi byta plats ?
kan du svara på det ?
kan du komma närmare ?
kan du komma närmre ?
kan ni komma närmare ?
kan ni komma närmre ?
kan du kontakta Tom ?
kan du beskriva den ?
kan du göra vad som helst ?
kan du förklara varför ?
kan du hantera det ?
kan du spela gitarr ?
kan du läsa arabiska ?
kan du reparera den här ?
kan du reparera det här ?
kan ni reparera det här ?
kan ni reparera den här ?
kan ni reparera denna ?
kan du reparera denna ?
kan du reparera detta ?
kan du säga det igen ?
kan du börja idag ?
kan du köra ännu ?
kan du över huvud taget simma ?
kom tillbaks om en vecka .
kom tillbaka om en vecka .
kom och träffa allihop .
kom till mötet .
kom på mötet .
kan jag tala med dig ?
kan du vara snäll och gå ?
kan du stanna bilen ?
kan du skriva under det här ?
kan du sakta ner ?
dela ut korten , Tom .
Förstör det här templet .
väckte jag er ?
gjorde Tom någonting ?
har Tom gjort någonting ?
köpte Tom den ?
har någon ringt mig ?
berättade någon för Tom ?
störtade planet ?
trodde du på Tom ?
tog du med frallor ?
gjorde du någonting ?
har ni gift er ?
gifte ni er ?
hade du drömmar ?
gav du dricks ?
har du gått ned i vikt ?
målade du de här ?
såg du någon ?
måste jag gå nu ?
får jag ändå betalt ?
gå inte nära dem .
har vi något val ?
behöver vi en plan B ?
tror du på det här ?
njuter du av att förlora ?
ger du lektioner ?
har du feber ?
har du något hus ?
har ni något hus ?
har du ett motto ?
har du en telefon ?
har ni en telefon ?
tycker du om att tälta ?
tycker du om löpning ?
tycker du om att springa ?
tycker du om hjortkött ?
tycker du om att promenera ?
känner du igen mig ?
ser du någonting ?
reser du ofta ?
tror Tom på mig ?
äter Tom vindruvor ?
ler Tom någonsin ?
har Tom kabel @-@ tv ?
ser Tom arg ut ?
ser Tom upprörd ut ?
simmar Tom ofta ?
spelar det någon roll ?
gör det verkligen ont ?
fungerar det ens ?
känns det där bra ?
skrämmer det dig ?
verkar det klokt ?
har du ont i huvudet ?
jobbar din fru ?
spela inte förvånad .
var inte så självisk .
gör inte så mot mig .
tappa inte den där koppen .
bli inte arg på mig .
bli inte arg på oss .
kom inte för nära .
tappa inte tilltron till mig .
avbryt inte Tom .
prata inte strunt .
rita en liten cirkel .
drick ditt te , Tom .
släpp kniven , Tom .
ät mer grönsaker .
alla sittplatser var upptagna .
alla applåderade .
alla ler .
alla är oroliga .
alla har ett namn .
alla skrattar .
alla står .
alla står upp .
allt är bättre .
allt är förstört .
Starta motorerna .
fixa en biljett åt mig .
kom bort därifrån .
gå bort därifrån .
kom tillbaks in i bilen .
kom tillbaks in i skåpbilen .
klä på dig fort .
klä på er fort .
Kläd på er fort .
Kläd på dig fort .
klä på dig snabbt .
klä på er snabbt .
Försvinn , ditt äckel .
ring efter en ambulans åt mig .
Försvinn från mina ägor .
skynda på , Tom .
Raska på , Tom .
ge Tom lite pengar .
ge Tom lite plats .
ge mig en till .
ge mig den där flaskan .
ge mig det där vapnet .
ge mig biljetterna .
ge mig tre timmar .
ge mig tre veckor .
ge mig din plånbok .
ge mig ditt vapen .
ge dem mitt nummer .
ge oss detaljerna .
gå och sök efter Tom .
gå och gör läxorna .
drick inte för mycket vin .
gå och hämta en tröja åt mig .
drick det nu , Tom .
gå på offensiven .
gissa hur lång jag är .
har Tom märkt någonting ännu ?
har den skadats ?
har jag blivit galen ?
har de gjort det ?
har du tolkat den ?
har du dechiffrerat den ?
har du provat det här ?
har du smakat det här ?
han säger alltid sådär .
han vände bort blicken .
han slog rekordet .
han brast i gråt .
han kan hjälpa dig .
han förnekade den uppgiften .
han kör en Ferrari .
han stiger upp klockan sju .
han steg på tåget .
han har ett gott hjärta .
han har gått för långt .
han har polisonger .
han låg på rygg .
han behöver de där pengarna .
han ljuger aldrig .
han kommer ofta sent .
han motsatte sig planen .
han festar för mycket .
han nådde sitt mål .
han gick i pension vid sextio .
han springer snabbast .
han satt i stolen .
han rakar sig varje dag .
han började svära .
han slutade plötsligt .
han stannade till plötsligt .
han kommer tillbaka sex .
han är lika stor som jag .
han är i femtioårsåldern .
hjälp mig att klä på mig .
hennes tal tråkade ut mig .
det är såhär vi gör .
du , jag har en idé .
du , kolla in det här .
du där , kom tillbaka .
hej , du ser jättebra ut .
hans biceps är jättestora .
hans idéer är galna .
jag kan inte komma på vad han heter .
håll i era hattar .
håll ut dina händer .
håll huvudet högt .
Älskling , är du skadad ?
det är kanske bättre att jag gör det .
ska vi tävla ?
det är ju hur bra som helst !
hur illa kan det vara ?
hur svårt skadad är Tom ?
hur ont gör det ?
hur kan jag nå Tom ?
hur ska jag kunna lita på dig ?
hur kan Tom göra så ?
hur kan Tom göra såhär ?
hur kan vi hjälpa Tom ?
hur kan vi hjälpa dig ?
hur kan vi stå till tjänst ?
hur kan vi bevisa det ?
hur kan vi rädda Tom ?
hur kan du vara säker ?
hur kan du göra sådär ?
hur kan du göra såhär ?
hur kan du hjälpa mig ?
hur skulle jag kunna göra det ?
hur djupt är det här ?
hur kunde jag missa det där ?
hur kunde jag missa det här ?
hur gjorde Tom det där ?
hur gjorde Tom det här ?
hur hittade Tom oss ?
vad tyckte Tom om den ?
hur tog Tom det ?
hur kom den hit ?
hur hände det där ?
hur hittade ni oss ?
hur hittade du oss ?
hur fick du slut på det ?
hur stoppade du det ?
hur överlevde du ?
Hurdan var din dag ?
hur ska jag förklara det ?
hur når jag NHK ?
hur gör de det ?
hur vet vi det ?
hur ska vi stoppa dem ?
hur lagar man den här ?
hur känner du Tom ?
hur känner ni Tom ?
hur säger man det ?
hur hjälper det oss ?
hur effektiv är den ?
hur långt borta är Tom ?
hur långt kom Tom ?
hur varmt blir det ?
på vilket sätt är det annorlunda ?
hur stora var de ?
hur länge har vi på oss ?
hur lång tid har vi ?
hur mycket förlorade jag ?
hur mycket äter du ?
hur mycket blir det ?
hur gammal är du nu ?
hur gammal är din son ?
hur var återträffen ?
hur var seminariet ?
hur ska du fly ?
hur ska du klara dig ?
hur ska ni klara er ?
hur skulle det hjälpa ?
hur skulle det se ut ?
hur skulle du reagera ?
jag beundrar ditt mod .
jag ringde nästan till Tom .
jag blev nästan rånad .
jag dödade nästan Tom .
jag var nära att döda Tom .
jag kysste nästan Tom .
det vet jag redan .
jag ångrar det redan .
jag sålde den där redan .
jag tar alltid bussen .
jag antecknar alltid .
så har jag alltid tyckt .
jag är också lärare .
jag är förföljd .
jag är inte din fiende .
jag är inte er fiende .
jag spelar gitarr .
jag är dålig på tennis .
jag skriver ett sms .
jag ber om ursäkt för Tom .
jag bad Tom att sluta .
jag vann över honom på schack .
jag slog honom på schack .
jag tror att Tom vet .
jag tror på hennes berättelse .
jag tror på mig själv .
jag köpte en sandwich .
jag köpte en dubbelmacka .
jag köpte lite grejer .
jag gjorde slut med Tom .
jag tog med mig lite vin .
jag tog med lunch till dig .
jag byggde ett nytt hus .
jag ringde polisen .
jag kom tillbaka för din skull .
jag kom för att säga hej .
jag kan komma klockan tre .
jag kan göra det åt dig .
jag kan göra det för dig .
jag kan stå upp för mig själv .
jag kan höra vinden .
jag kan hålla en hemlighet .
jag kan åka med Tom .
jag kan stoppa läckan .
jag känner doften av blommor .
det doftar blommor .
jag kan ännu göra det .
jag kan överleva ensam .
jag kan föra hem Tom .
jag kan förstå det .
jag kan vänta här ute .
jag kan inte svara på det .
jag kan inte ändra på det .
jag kan inte kontakta Tom .
jag får inte kontakt med Tom .
jag kan inte få kontakt med Tom .
jag kan inte kontrollera Tom .
jag kan inte göra mer .
jag kan inte göra det själv .
jag klarar det inte själv .
jag kan inte göra det i dag .
jag klarar det inte i dag .
jag klara det inte nu .
jag kan inte rita en fågel .
jag kan inte gå tillbaka nu .
jag kan inte titta på Tom .
jag klarar inte av lögnare .
jag står inte ut med lögnare .
jag kollade måttet .
jag kan ha tagit fel .
jag kan ha fel .
jag kunde göra det igen .
jag kunde äta en häst .
jag kan komma med dig .
jag kunde knappt vänta .
jag kan förlora mitt jobb .
jag kan tala med Tom .
jag skulle kunna tala med Tom .
jag grät hela morgonen .
jag inredde mitt rum .
jag kollade upp några saker .
jag forskade lite .
det gjorde jag för länge sedan .
jag gjorde det en gång .
jag behövde inte gå .
jag behövde inte åka .
jag var inte tvungen att gå .
jag var inte tvungen att åka .
jag sov inte bra .
jag håller inte med Tom .
jag håller inte med dig .
jag behöver en tjänst .
jag behöver verkligen din hjälp .
jag förstår inte .
jag ber faktiskt ibland .
jag litar verkligen på dig , Tom .
jag oroar mig verkligen för det .
jag går inte ut så ofta .
jag har inte ett öre .
jag har ingen kostym .
jag vet egentligen inte .
jag vet inte riktigt .
jag äter mycket kött .
jag äter med händerna .
jag tyckte om den här boken .
jag känner mig tom inombords .
jag känner mig liksom lite sjuk .
jag känner mig som en slav .
jag känner för att vänta .
jag känner mig väldigt olycklig .
jag fixar trasiga radioapparater .
jag följde efter Tom hit .
jag bar mig ohyfsat åt .
jag glömde att fråga Tom .
jag gav Tom ett äpple .
jag fattar vad du menar .
jag har gift mig igen .
jag gifte mig ung .
jag blev riktigt hungrig .
jag fick den av Tom .
jag köpte någonting åt dig .
jag har köpt någonting åt dig .
jag åt en hyfsad måltid .
jag kände på mig det .
jag hade en förkänsla av det .
jag hade mina misstankar .
jag hade ett sista hopp .
jag var tvungen att göra min plikt .
jag var tvungen att hyra en bil .
jag hatar väckarklockor .
jag hatar att vara chef .
jag hatar att vara singel .
jag hatar att vara dum .
jag hatar det där så mycket .
jag hatar den där trumpeten .
jag hatar det här vädret .
jag hatar de där sakerna .
jag hatar de där .
jag hatade det först .
jag har en stor familj .
jag har ett handikapp .
jag har en flickvän .
jag har en jättebra idé .
jag har ett ledigt rum .
jag har styv nacke .
jag har ett öppet sinne .
jag har en annan idé .
jag har en annan plan .
jag har varit i Rom .
jag har räkningar att betala .
jag har klardrömmar .
jag har ett eget hus .
jag har ingenting att invända .
jag har ingenting annat .
jag har en sådan .
jag har en fråga .
jag har bara en penna .
jag har flera kepsar .
jag har ett flertal kepsar .
jag har tennisarmbåge .
jag måste ändra den .
jag måste göra det nu .
jag måste göra mitt jobb .
jag måste ge mig i väg .
jag måste gå och byta om .
jag måste gå och byta kläder .
jag måste gå nu .
jag måste bege mig nu .
jag måste ge mig av nu .
jag måste lämna dig .
jag måste sjappa .
jag måste ge mig av .
jag måste sluta upp med det här .
jag måste få ett slut på det här .
jag måste studera nu .
jag måste plugga nu .
jag måste lita på Tom .
jag har dig att tacka .
jag har era biljetter .
jag hörde att det var trevligt .
jag hörde meddelandet .
jag gömde mig under sängen .
jag hoppas att Tom hjälper mig .
jag hoppas att Tom har fel .
jag hoppas att Tom säger ja .
jag hoppas att det ordnar sig .
jag hoppas att de gillar mig .
jag hoppas att du kan hjälpa till .
jag hoppas att du hittar Tom .
jag hoppas att du tycker om Tom .
jag hoppas att du har rätt .
jag gjorde mig illa idag .
jag har för avsikt att göra det .
jag rengjorde den här nyss .
jag klippte nyss naglarna .
jag bara älskar blommor .
jag vill bara ha svar .
jag vill bara veta .
jag vill bara prata .
det visste jag redan .
jag visste att du skulle bli arg .
jag vet att Tom har rätt .
det vet jag redan .
jag vet vad de är för ena .
jag känner de här personerna .
jag vet att det här är svårt .
jag vet att detta är svårt .
jag vet att det är svårt .
jag vet vad som är rätt .
jag vet var hon är .
jag vet att du mår dåligt .
jag vet att du har rätt .
jag vet att du är upprörd .
jag vet att ni är upprörda .
jag känner er bror .
jag tycker om fattiga riddare .
jag gillar dina speglar .
jag gillade ditt tal .
jag älskar kinamat .
jag älskar kinesisk mat .
jag älskar det programmet .
jag älskar det här företaget .
jag älskar den här bilden .
jag tjänar 100 euro om dagen .
jag träffade honom i går .
jag kanske kommer att prata med Tom .
jag kanske pratar med Tom .
jag måste bege mig nu .
jag måste ge mig av nu .
jag måste gå nu .
jag måste göra någonting .
jag måste åka någonstans .
jag måste lära mig franska .
jag måste jobba ikväll .
jag behöver en ordbok .
jag behöver en flickvän .
jag behöver en stor tjänst .
jag behöver hjälp här inne .
jag behöver svar .
jag behöver bilnycklarna .
jag behöver lösenordet .
jag måste komma hem .
jag måste få en penna .
jag behöver dig en sekund .
du måste köra .
du måste gå .
jag kunde aldrig göra det .
jag tvivlade aldrig på dig .
jag ljög aldrig för Tom .
jag börjar aldrig slåss .
jag rörde aldrig Tom .
jag ville aldrig ha den här .
jag önskar bara hjälpa .
jag vill bara vara till hjälp .
jag polerade mina skor .
jag låtsades arbeta .
jag ringde på dörrklockan .
jag har verkligen otur !
det tvivlar jag faktiskt på .
jag kommer ihåg allt det där .
jag minns allt det där .
jag kommer ihåg den här kartan .
jag omarbetade min teori .
jag reviderade min teori .
jag sa god morgon .
god morgon , sa jag .
jag såg henne i går .
jag såg en igår .
jag såg ett igår .
jag såg vad som hände .
jag träffar Tom varje dag .
jag ser Tom varje dag .
jag borde vila .
jag borde inte vara här .
jag pratar franska också .
jag stal den från Tom .
jag stal det från Tom .
jag studerar konsthistoria .
jag kände mig plötsligt gammal .
jag föreslår att du skyndar dig .
jag lärde Tom franska .
jag tror att jag satt på den .
jag tror att jag satte mig på den .
jag tror att jag är förälskad .
jag tror att jag är kär .
jag tycker att du är trevlig .
jag tycker att du är snäll .
jag tänkte på Tom .
jag trodde att vi hade kommit överens .
jag sa åt Tom att ta det lugnt .
jag sa åt dig att gå .
jag sa åt er att gå .
jag sa åt dig att ge dig iväg .
jag sa åt er att ge er iväg .
jag tog den här bilden .
jag ansträngde mig verkligen .
jag försökte varna dig .
jag försökte varna er .
jag litar på läraren .
jag vill ha en glass .
jag vill be om ursäkt .
jag vill komma hem .
jag vill äta pizza .
jag vill gifta mig med henne .
jag vill att du dansar .
jag var självisk .
jag följde efter dig .
jag var på dåligt humör .
jag gissade bara .
jag fick en judisk uppfostran .
jag var jättehungrig .
jag tog ett bad .
jag tvättade min T @-@ shirt .
jag diskade .
jag tvättade lakanen .
jag var inte ens där .
jag såg Tom ge sig av .
jag gick tillbaka till jobbet .
jag kommer tillbaka snart .
jag går om du går .
jag önskar att jag hade ett band .
jag önskar att jag hade en tvilling .
jag önskar att jag förstod .
jag önskar att Tom var här .
jag önskar att Tom vore här .
jag skrev det brevet .
det skulle gå bra för mig .
jag hjälper gärna till .
jag skulle dö utan dig .
jag skulle dö utan er .
jag skulle vilja träffa Tom .
jag skulle vilja se Tom .
jag ska vara snäll mot Tom .
jag åker gärna .
jag kommer att vara utanför stan .
jag ska köpa en öl till Tom .
jag ringer efter en taxi åt dig .
jag ringer en taxi åt dig .
jag gör som jag vill .
jag ska göra som du önskar .
jag gör som jag vill .
jag hämtar den åt dig .
jag hämtar läkaren .
jag hämtar stegen .
jag hämtar de andra .
jag vänjer mig .
jag ska hämta en öl åt dig .
jag ska ge dem tillbaka .
jag ska gå och hämta Tom .
jag går och byter om .
jag går om en minut .
jag tar dina väskor .
jag vaktar dörren .
jag kommer att sakna dig mycket .
jag betalar på mitt eget sätt .
jag berättar för Tom senare .
jag ska berätta för Tom senare .
jag är lite hungrig .
jag är socialarbetare .
jag är socialvårdare .
jag är en främling här .
jag är helt säker !
jag är oskyldig .
jag är på en servicestation för lastbilar .
jag blir hämtad .
jag blir upphämtad .
jag blir uppraggad .
jag håller på att bli uppraggad .
jag gör det själv .
jag dricker kaffe .
jag är glad att kunna hjälpa till .
jag är glad att vi såg Tom .
jag åker in till stan .
jag ska börja banta .
jag ska laga den .
jag ska gå nu .
jag kommer att gå nu .
jag går nu .
jag är på väg åt det hållet .
jag är något av en ensamvarg .
jag är inte bra för dig .
jag är ingen konstkännare .
jag är inte ett dugg trött .
jag är inte bra på att ljuga .
jag är inte alls upptagen .
jag är inte alls frisk .
jag är inte elak .
jag kommer inte att gå .
jag har inte ont .
jag har inte ont någonstans .
jag är inte stolt över det .
jag är inte så säker nu .
jag är på väg dit .
jag är bara en kund .
jag är så stolt över dig .
jag är din nya advokat .
jag har lånat en bil .
jag har några till .
jag har en fråga .
jag har jättegoda nyheter .
jag har fått lite idéer .
jag har tre barn .
jag måste vara fri .
jag måste återvända .
jag måste gå tillbaka .
jag måste gå , Tom .
jag har jobb att sköta .
jag har haft en dålig vecka .
jag har precis kommit hem .
jag har precis ätit lunch .
jag har nyss ätit lunch .
är Tom fortfarande singel ?
är någonting av detta verkligt ?
är någonting av detta sant ?
är allt där ?
är det ett ja eller ett nej ?
är vädret fint ?
är den här radion din ?
är detta äkta silver ?
är inte det planen ?
är det inte det som är planen ?
det stör mig mycket .
det kostade mig skjortan .
det kan vara ett påhitt .
det hände så fort .
det hände så snabbt .
det är iskallt .
det kommer att komma snö .
det kommer att snöa .
det måste bli gjort .
det regnade i går .
det tog hela kvällen .
det var nästan roligt .
det var ganska roligt .
det var riktigt roligt .
det var oförlåtligt .
jag höll på i flera dagar .
det blir en lång dag .
det är en av livets realiteter .
det är en enda röra här inne .
den är ungefär så här stor .
det hela är ett stort skämt .
det hela är nytt för mig .
klockan är redan elva .
det är svårt att acceptera .
det är svårt att motstå .
det är min gåva till dig .
det är ingen dålig affär .
det är ingen dålig idé .
det är ingen dålig plan .
det är inte bara en penna .
det är en del av mitt arbete .
det är kvavt här inne .
det är kvalmigt här inne .
det är dags att gå nu .
det är väldigt varmt idag .
det är väldigt varmt i dag .
Jesus svarade dem .
berätta bara inte för Tom .
följ bara mitt exempel .
kom in och sätt dig i bilen bara .
sätt dig i bilen bara .
sätt igång nu bara .
ge den åt Tom bara .
ge mig ett handtag bara .
ge mig min pistol bara .
gå och lägg dig igen nu .
håll ett öga på dem .
det får räcka för i dag .
ska vi sätta punkt här .
kom så går vi upp på däck .
låt Tom prata .
vi pratar engelska .
se på vad jag har lagat .
se vad jag har köpt åt dig .
många människor gör detta .
kan jag ringa upp dig senare ?
jag kanske somnade .
Apor klättrar i träd .
mer kaffe , tack .
kan jag få mer kaffe ?
min katt älskar räkor .
min pappa tycker om tennis .
det ringer i mina öron .
mina fingrar är domnade .
mina fingrar har domnat .
mitt hår är så smutsigt !
mitt hår är för långt .
mina händer är kladdiga .
mitt hus är hemsökt .
det spökar i mitt hus .
jag heter också Tom .
mina nya skor knarrar .
min brorsdotter är sjuksköterska .
min systerdotter är sjuksköterska .
mitt te är för sött .
mina lärare tycker om mig .
min dragkedja fastnade .
nästa person , tack !
ingen kom med mig .
ingen har någonting .
ingen tycker om att förlora .
ingen bryr sig egentligen .
det är ingen som faktiskt vet .
ingen kommer att bli skadad .
ingen kommer att överleva .
ingen hackade på mig .
ingen väntar på mig .
ingen skulle se oss .
det var ingen som ville ta emot oss .
ingen skriver till mig .
ingenting av det var verkligt .
ingenting av det var äkta .
ingenting kan stoppa den .
ingenting kan stoppa oss .
det är ingenting på gång .
nu kan jag dö lycklig .
jag känner mig lättad nu .
kom hit nu .
öppna dina ögon nu .
en av oss kunde vinna .
en av oss skulle kunna vinna .
en av er ljuger .
folk älskar frihet .
gör det för mig är du snäll .
var snäll och tala långsamt .
ta på dig en fin klänning .
vila dig här en stund .
Vässa din penna .
hon har inte råd med det .
hon gjorde rätt bra ifrån sig .
hon har gått och lagt sig .
hon har vackra ögon .
hon har mässlingen .
hon är mörkhyad .
hon fortsatte prata .
hon går sällan ut .
hon älskar honom fortfarande .
hon är en drama queen .
så vad ska jag göra nu ?
någon satte dit honom .
förr eller senare kommer vi att veta .
stanna där du är !
stanna där ni är !
sluta kalla mig för Tom .
sluta anmärka på Tom .
sluta hacka på Tom .
ta några dagar ledigt .
ta av dig skorna .
ta av er skorna .
säg till Tom att jag älskar honom .
berätta för Tom att jag älskar honom .
berätta sanningen för dem .
tack för informationen .
det låter logiskt .
det var en bra dag .
det är okej med mig .
det var så jag gjorde det .
det är så jag ser det .
det är så vi gör det .
det är så vi brukar göra .
bussen blir kanske sen .
hunden åt upp min sko .
hunden följde efter mig .
hunden blöder .
slutet är i sikte .
garaget är dammigt .
flickan hoppar .
huset är jättestökigt .
tanken är inte ny .
idén är inte ny .
sjön låg frusen .
sjön var tillfrusen .
orsaken är klar .
skeppet sjunker .
strumporna luktar illa .
Utsikten är fantastisk .
terapi fungerade inte .
det måste finnas ett sätt .
det finns ett villkor .
det finns ingen hiss .
dessa är reglerna .
de är kristna .
de tror på Gud .
de kan inte stoppa oss .
de såg förskräckta ut .
de började skjuta .
de kommer över det .
de kommer nog över det .
saker har förändrats .
det här är ett stort hus .
det här är lite läskigt .
det här är en guldgruva .
det här är en bra föreställning .
det här är en bra show .
det här är en bra plats .
det här är en lång lista .
det här är en trevlig plats .
det här är ett sjukt skämt .
det här är en gammal regel .
det här är lätt för mig .
det här är fantastiskt .
detta är deras hus .
det här är deras hus .
det här är väldigt läskigt .
det här måste vara ett skämt .
den här är speciell .
det här borde vara enkelt .
den här duger fint .
det är mina order .
det där är mina saker .
det är riskerna .
det är reglerna .
sådana är reglerna .
tiden verkade stanna .
Tom hade med sig blommor .
Tom kan köra bil .
Tom skrämde mig inte .
Tom äter som en gris .
Tom blev generad .
Tom högg tag i sin väska .
Tom grep tag i sin väska .
Tom ryckte till sig sin väska .
Tom hade en mardröm .
Tom hade mycket att göra .
Tom hörde fotsteg .
Tom höll Mary tätt .
Tom hjälpte oss mycket .
Tom la på i örat på Mary .
Tom lade på i örat på Mary .
Tom skadade sig .
Tom är en smart kille .
Tom är lite udda .
Tom äter långsamt .
Tom är tillgiven .
Tom är kärleksfull .
Tom är redan hemma .
Tom är tillbaka i stan .
Tom är grälsjuk .
Tom är besviken .
Tom är missnöjd .
Tom är missbelåten .
Tom ignorerar dig .
Tom är uppe på vinden .
Tom ligger i sängen .
Tom är flerspråkig .
Tom är verkligen ledsen .
Tom är högerhänt .
Tom sover fortfarande .
Tom gråter fortfarande .
Tom är fortfarande singel .
Tom är deras ledare .
Tom är för långt borta .
Tom är ingen turist .
Tom är inte turist .
Tom andas inte .
det är inte Tom som bestämmer .
Tom behöll min tändare .
Tom gick vidare .
Tom fortsatte gå .
Tom skrattade åt Mary .
Tom gillade den idén .
Tom tyckte om den idén .
Tom tycker om spagetti .
Tom gillar spagetti .
Tom tycker om att resa .
Tom bor på en båt .
Tom såg skräckslagen ut .
Tom ser lättad ut .
Tom ser annorlunda ut .
Tom ser äcklad ut .
Tom ser utmattad ut .
Tom ser utpumpad ut .
Tom ser slut ut .
Tom tog ett beslut .
Tom fattade ett beslut .
Tom valde .
Tom gjorde sitt val .
Tom fick mig att göra det .
Tom måste stoppas .
Tom behövde pengar .
Tom behövde kontanter .
Tom kom aldrig tillbaka .
Tom nickade tyst .
Tom öppnade dörren .
Tom äger den här bostaden .
Tom vägrar att prata .
Tom rullade med ögonen .
Tom himlade med ögonen .
Tom satt på trottoarkanten .
Tom sade åt oss att vänta .
Tom blev avvisad .
Tom fick avslag .
Tom fick nej .
Tom fick korgen .
Tom är en sympatisk kille .
sänk volymen på radion .
vänta i bilen , okej ?
vi har alla ett pris .
vi äter lunch .
vi kan ta itu med det .
vi kan skaffa hjälp åt dig .
vi kan hjälpa Tom nu .
vi kan få det att fungera .
vi kunde behöva lite hjälp .
vi gjorde det i skolan .
vi skrev faktiskt till dig .
vi har ingen bil .
vi har ingen katt .
vi har ingen hund .
vi kom hit i tid .
vi hann hit i tid .
vi hamnade i bråk .
vi åt en stor middag .
vi hade ett stort gräl .
vi hade jätteroligt .
vi har ett jobb att göra .
vi måste ringa Tom .
vi måste ta reda på .
vi måste få reda på det .
du måste flytta på dig nu .
du måste flytta nu .
vi måste stoppa Tom .
vi måste berätta för Tom .
vi måste berätta det för Tom .
vi måste prova det här .
vi måste jobba nu .
vi måste arbeta nu .
vi vet vem du är .
vi älskar dig så mycket .
vi måste göra det igen .
vi måste gå .
vi måste komma bort .
vi måste få hjälp .
vi måste hjälpa Tom .
vi måste stoppa Tom .
vi måste jobba nu .
vi borde sätta igång .
vi borde komma igång .
vi borde ge oss av .
vi reste till fots .
vi var nästan färdiga .
vi var nästan klara .
vi var i parken .
vi var vid parken .
vi var på parkeringen .
vi skojade bara .
vi var väldigt hungriga .
vi ska nog gå nu .
vi ska göra allt vi kan .
vi ska göra som du säger .
vi ska göra oss av med den .
vi hämtar lite till .
vi ska göra ett försök .
vi håller kontakt .
vi är båda studenter .
vi går ut nu .
vi måste åka nu .
vi måste prova det .
vilken fantastisk middag !
vilken hemsk dag !
vad har jag för alternativ ?
vad har de på gång ?
vad äter du ?
vad ska du ta ?
vad har du för planer ?
Vilka är dina villkor ?
vad hände med dem ?
vad kan jag säga till Tom ?
vad kan du göra nu ?
vilken färg är de ?
vad kan Tom mena ?
vad kunde vara fel ?
vad förväntade sig Tom ?
vad hade Tom förväntat sig ?
vad glömde Tom ?
vad köpte Tom till mig ?
vad slog han upp ?
vad bevisade det ?
vad erbjöd de ?
vad hade de att erbjuda ?
vad svarade de ?
vad tyckte de ?
hur ser jag ut ?
vad ska jag säga först ?
vad ska vi göra först ?
vad säger vi till Tom ?
vad tror du på ?
vad jobbar ni med ?
vad är du skyldig Tom ?
vad ser du nu ?
vad föreslår du ?
vad undervisar Tom i ?
vad lär Tom ut ?
vad anser Tom ?
vad tycker Tom ?
vad spelar det för roll ?
vad kostar det ?
vad mer kan jag säga ?
vad annat gör du ?
vad annat behövs ?
vad hände med den ?
vad har du hört ?
vad har du tagit ?
vad gör vi om Tom säger nej ?
vad har hon för problem ?
vad är det med henne ?
vad har han för problem ?
vad är det med honom ?
vad finns i den här lådan ?
vad har vi för problem ?
vad är populärt nu ?
vad är inne nu ?
vad är på modet nu ?
vad är ditt val ?
vilken har du valt ?
vilken väljer du ?
Vilka vackra blommor !
vad mer kan jag be om ?
vad mer kan jag säga ?
vad mer kan vi göra ?
Vilka fina blommor !
vad var Toms plan ?
vad hade du på gång ?
vad är du bra på ?
gjort är gjort .
vad är det som händer nu ?
vad har tagit åt dig ?
vad är ditt problem ?
när kan vi flytta in ?
när kan vi träffa Tom ?
när rymde Tom ?
när får vi betalt ?
när ska Tom vara tillbaka ?
var är mina saker ?
var är våra sittplatser ?
vart ska du ta vägen ?
var är du i dag ?
var är era barn ?
var kan jag hitta den ?
var kan jag tvätta mig ?
var gjorde du det ?
var använder man den ?
vart är smöret ?
var ligger museet ?
var ligger toaletten ?
var ligger ditt hus ?
var ska vi träffas ?
var är min golfbag ?
var ligger flygplatsen ?
var är din jacka ?
vilket lag kommer att vinna ?
vem kan hindra oss nu ?
vem är din lärare ?
vem brukade göra detta ?
vem brukade göra det här ?
vems glas är det här ?
vems idé var det ?
vems telefon är det där ?
vems skjorta är det här ?
varför är jag fortfarande här ?
varför är du hemma ?
varför är ni hemma ?
varför är du i stan ?
vad skakar du för ?
varför skakar du ?
varför skakar ni ?
varför är du så säker ?
varför är du med mig ?
varför ta upp det nu ?
varför kysste Tom mig ?
varför sa vi det där ?
varför sa vi sådär ?
varför gav du upp ?
varför gick du din väg ?
varför åkte du iväg ?
varför hjälpte du mig ?
varför valde du mig ?
varför sa du ja ?
varför sålde du den ?
varför kom du förbi ?
varför måste jag gå ?
varför gör de så ?
varför frågar du det ?
varför undrar du ?
varför hatar ni Tom ?
varför tycker du om Tom ?
varför åker inte Tom ?
varför ger sig Tom inte iväg ?
skulle Tom gilla det ?
skulle Tom tycka om det ?
du är i otakt .
du kan lita på Tom .
du kan tala med Tom .
du kan inte neka det .
du gjorde ett jättebra jobb .
du ger mig så mycket .
ni måste gå .
du hatar Tom , eller hur ?
ni hatar Tom , eller hur ?
du har ett bra arbete .
du måste hålla ut .
du måste berätta för oss .
du måste berätta det för oss .
du har jobb att göra .
du ser blek ut idag .
du måste gå tillbaka .
du måste återvända .
du måste gå hem .
du måste hålla tyst .
du var en duktig pojke .
ni kommer att behöva en nyckel .
du skulle vara bra på det .
du kommer att avslöja mig .
du är så vacker .
ni är så vackra .
du är en sådan flörtis .
du är anhållen .
du har ätit tillräckligt .
ni har ätit tillräckligt .
du har en timme på dig .
din bil brinner .
du är fin i håret .
era skor är här .
en kopp te , tack .
pianon är dyra .
det är dyrt med pianon .
alla mina saker är här .
alla mina grejer är här .
alla mina grejor är här .
allting måste förgå .
alla tre män log .
är jag misstänkt ?
vad som helst är möjligt .
Apor är intelligenta .
är det där mina glasögon ?
ska vi sätta igång snart ?
ska vi börja snart ?
är du rädd för mig ?
är du färdig ännu ?
följer ni efter mig ?
håller du på bli tokig ?
fattar du det här ?
tänker du åka snart ?
har ni öppet ikväll ?
är du pensionerad , Tom ?
tänker du stanna kvar , Tom ?
är du deras mamma ?
är du olycklig , Tom ?
ska du gå hem ?
jobbar du hårt ?
var tysta båda två .
hämta mig en torr handduk .
hämta hit de där männen .
får jag fråga vad det är ?
får jag bjuda dig på middag ?
kan jag ringa upp dig ?
kan jag köra dig hem ?
kan jag träffa dig där ?
får jag se rapporten ?
får jag se dina händer ?
kan jag börja imorgon ?
kan jag tänka på det ?
kan jag tänka på saken ?
kan folk köpa de här ?
har vi råd med det nu ?
kan vi gå och ta en promenad ?
kan vi intervjua Tom ?
kan du beskriva honom ?
kan du göra det åt mig ?
kan du göra det för mig ?
kan du laga en toalett ?
klarar du dig på egen hand ?
kan du översätta det ?
kan vi inte göra något ?
kan vi inte göra någonting ?
vi ses senare , Tom .
vi hörs senare , Tom .
blunda , Tom .
Kyla gör armar och ben stela .
kom och hjälp mig .
kom och hälsa på mig snart .
kom och ta en titt .
kom tillbaks om en timme .
kom tillbaka om en timme .
kom hit , unge man .
kom in en minut .
kom ut därifrån nu .
var snäll och kom med oss .
Bomull absorberar vatten .
kunde jag få låna en såg ?
missade jag någonting ?
gjorde jag faktiskt det ?
gjorde Tom sig illa ?
berättade Tom för någon ?
Hotade Tom dig ?
gjorde någon sig illa ?
fick han ett kvitto ?
gick det bra i dag ?
slog någon Tom ?
körde vi på någonting ?
åt du något ?
frågade du ut Tom ?
Hotade du Tom ?
vann du kapplöpningen ?
vann du kappkörningen ?
visste du inte det ?
måste jag göra det ?
måste jag betala er ?
behöver jag betala dig ?
behöver jag betala er ?
gör det någon annanstans .
gör inte andra illa .
har de vapen ?
har vi en försäkring ?
bär du på vapen ?
har du lust med det ?
har du någon familj ?
har ni någon familj ?
har du ett garage ?
har du några kontanter ?
har du något käk ?
har du läxor ?
har du några skador ?
har du boken ?
tycker du om rödvin ?
tycker du om att studera ?
tycker du om ditt jobb ?
trivs du på ditt jobb ?
Mediterar du , Tom ?
går det bra att jag sitter ?
behöver du någonting ?
behöver ni någonting ?
äger du ett handeldvapen ?
äger du ett eldhandvapen ?
känner du igen honom ?
kommer du ihåg det ?
minns du dem ?
kommer du ihåg dem ?
förstår du mig ?
vill ni ha en banan ?
vill ni ha ett äpple ?
arbetar ni tillsammans ?
överraskar det dig ?
låter det vettigt ?
fungerar den här ännu ?
fungerar den här ?
fungerar den här apparaten ?
var inte så dramatisk .
var inte så negativa .
var inte en sådan barnunge .
glöm inte att rösta .
lämna mig inte ensam .
låt inte tom skrika .
rör inte mina grejor .
rör inte mina grejer .
rör inte mina prylar .
rör inte mina saker .
vill du inte åka ?
till och med mamma vet om det .
varje familj har en sådan .
alla gör det .
alla är här nu .
alla höll sig lugna .
Samtliga höll sig lugna .
alla sa nej till Tom .
allt gick bra .
allt har förändrats .
ursäkta mig ett ögonblick .
äntligen är det fredag .
äntligen fredag .
hitta någonstans att sitta .
fokusera på nuläget .
lämna min son i fred .
ta kontakt med mig .
gör dig färdig för skolan .
ge den en timme till .
ge mig en dag eller två .
ge mig en till spik .
ge mig lösenordet .
ge mig de där .
ge mig era plånböcker .
ge mig era vapen .
gå och fråga Tom .
prova den nu då .
gå och snygga till dig .
gå och fyll ispåsen .
gå och hämta ditt pass .
gå hem till din fru .
Fortsätt med ditt arbete .
Grabba tag i någonting .
ge mig de där pappren .
har Tom redan åkt ?
har Tom varit hjälpsam ?
har Tom blivit skadad ?
har Tom blivit nedsövd ?
har Tom slutat röka ?
har han pratat med dig ?
ta en drink med mig .
ha en trevlig dag , Tom .
har du förrått oss ?
har du svikit oss ?
har du förlåtit mig ?
har du gått ner i vikt ?
har du sett min son ?
har ni sett min son ?
har du börjat ännu ?
han spelar alltid bra .
han jobbar alltid hårt .
han bad om min hjälp .
han har byggt ett nytt hus .
han byggde ett nytt hus .
han hade femtio dollar .
han har hår på bröstet .
han har en stor lastbil .
han är en blid natur .
han är en god simmare .
han är på väg att gå .
han är alltid med mig .
han är sitt vanliga jag .
han är inte här längre .
han läser en bok .
han tycker mycket om musik .
han gillar den här gitarren .
han bor i Nagasaki .
han ser lite trött ut .
han berättade aldrig för någon .
han spelar ofta piano .
han rusade in i rummet .
han tog av sig skjortan .
han reparerade näten .
han pratade väldigt högt .
han jobbar på banken .
han har en vit katt .
han är på sjukhuset .
han är bara en amatör .
han är aldrig nöjd .
här är några idiomatiska uttryck .
här är ditt kvitto .
vänta en sekund .
skulle det smaka med en smörgås ?
hur har Tom och Mary det ?
hur svårt skadad var Tom ?
hur stort är ditt rum ?
hur kan jag hjälpa till ?
hur kan jag vara till hjälp ?
hur kan de göra så ?
hur kan detta vara sant ?
hur kan det vara sant ?
hur kan vi stoppa dem ?
hur kan vi tacka er ?
hur kan vi tacka dig ?
hur kan du äta det där ?
hur skulle jag kunna hata Tom ?
hur fick Tom reda på det ?
hur kom Tom hem ?
hur blev Tom skadad ?
hur blev Tom rik ?
hur knäckte du den ?
hur hade du sönder den ?
hur hittade du Tom ?
hur fick du reda på det ?
hur fick du tag i den här ?
hur gick det för dig ?
hur träffade du honom ?
hur gick träffen ?
hur gör föräldrar det ?
hur känner du dig , Tom ?
hur vet du det ?
hur gör Tom det där ?
hur långt skulle Tom gå ?
hur fort kan du springa ?
hur fort sprang Tom ?
hur snabbt sprang Tom ?
hur är detta relevant ?
hur lång tid har vi ?
hur lång tid har vi på oss ?
hur många fick du ?
hur många fick du tag på ?
hur många vill ni ha ?
hur mycket såg du ?
hur mycket vet du ?
hur mycket tjänar du ?
hur mycket vill ni ha ?
hur mycket kostar en biljett ?
vad kostar en öl ?
hur hög är hyran ?
hur mycket är för mycket ?
hur gamla är ni ?
hur gammal är du , Tom ?
hur gammal var Tom då ?
hur dödades de ?
hur är det med din fru , Tom ?
jag jobbar faktiskt här .
jag känner mig nästan skyldig .
jag tror på det redan .
jag ringde redan till Tom .
jag provade det där redan .
jag väntar på min tur .
jag skriver en roman .
jag anlände igår kväll .
jag anlände i går kväll .
jag bad Tom att gå .
jag bad om att få pengarna tillbaka .
jag besökte festen .
jag slår vad om att jag blir klar först .
den här ska nog fungera .
jag köpte någonting smått att äta åt dem .
jag hade sönder en vas idag .
jag tog med en present till dig .
jag brast ut i skratt .
jag kan äta den här inne .
jag kan knappt andas .
jag kan knappt se honom .
jag kan hjälpa med det där .
jag kan hjälpa till med det där .
jag klarar mig , tack .
jag kan ännu hjälpa dig .
jag kan skjutsa dig dit .
jag kan tala om det för dig senare .
jag kan förstå dig .
jag kan inte sjunga en ren ton .
jag kan inte komma i kväll .
jag kan inte bekräfta det .
jag kan inte övertyga Tom .
jag kan inte heller dansa .
jag kan inte dansa heller .
jag kan inte bli inblandad .
jag hör ingenting .
jag kan inte höra någonting .
jag kan inte leva med det .
jag kan inte riskera någonting .
jag kan inte ta några risker .
jag valde en annan väg .
jag valde en annan stig .
jag valde att inte åka .
jag kunde knappt prata .
jag kan vara misstänkt .
jag kan dö imorgon .
jag kan gå dit nu .
jag skulle kunna hjälpa dig .
jag kunde inte bry mig mindre .
jag skulle inte kunna bry mig mindre .
det rör mig inte i ryggen .
jag designade den själv .
jag hittade faktiskt någonting .
jag hittade faktiskt en sak .
jag gick inte och la mig .
jag gick inte med Tom .
jag följde inte med Tom .
jag dödade inte någon .
jag gör det hela tiden .
jag tror inte på det .
jag förtjänar inte detta .
jag förtjänar inte det här .
jag hör ingenting .
jag hör inte ett skvatt .
jag kan inte engelska .
jag har inget emot att hjälpa till .
jag känner inte igen det .
jag känner inte igen den .
jag litar inte på någon .
jag vill inte laga mat .
jag vill inte leva .
jag vill inte leka .
jag vill inte vila .
jag faxade en karta åt Tom .
jag känner mig lite öm .
jag känner mig säker på det .
jag känner mig väldigt förrådd .
jag tyckte synd om Tom .
jag följde efter Tom dit .
jag glömde att ringa Tom .
jag glömde att kolla på det .
jag går vart jag vill .
jag hämtade lite vatten åt Tom .
jag fick B i fysik .
jag fick C i engelska .
jag fick betalt igår .
jag fick lön igår .
jag steg upp tidigt idag .
jag antar att Tom har rätt .
jag antar att du har rätt .
jag hade en bra semester .
jag åt lunch med Tom .
vi var tvungna att fortsätta .
jag råkar gilla Tom .
jag hårdkokte ett ägg .
jag hårdkokade ett ägg .
jag går nästan aldrig ut .
jag hatar skräckfilmer .
jag avskyr skräckfilmer .
jag har en skuld att betala .
jag har några minuter .
jag har en hushållerska .
jag har hushållerska .
jag har ont i halsen .
jag har en inbjudan .
jag har ryggproblem .
jag har hemska nyheter .
jag har vänner där .
jag måste bege mig nu .
jag har massor av pengar .
jag har min egen teori .
jag har ingen statistik .
jag har så många idéer .
jag har sådan otur .
jag måste ge mig i väg .
jag måste gå och göra det här .
jag måste börja om .
jag måste jobba idag .
jag har två döttrar .
jag har vad du behöver .
jag har inte fått den än .
jag har hört att Tom hatar dig .
jag hörde att jag behövdes .
jag hörde vad som har hänt .
jag hörde de dåliga nyheterna .
jag hörde frågan .
jag hoppas att jag kan göra det här .
jag hoppas att de tyckte om mig .
jag hoppas att du tycker om den här .
jag hoppas att du är hungrig .
Inledningsvis hatade jag det .
jag skar mig just i fingret .
jag skar mig nyss i fingret .
jag fick just en vän .
jag behöver bara en minut .
jag visste att jag måste sluta .
jag visste att det inte var du .
jag visste att det inte var ni .
jag visste att du skulle vara upptagen .
jag visste att du skulle gilla det .
jag visste att du skulle gilla den .
jag visste att du skulle tycka om det .
jag visste att du skulle tycka om den .
jag visste att du skulle sakna mig .
jag visste att ni skulle sakna mig .
jag vet att jag kan göra mer .
jag vet allt om dig .
jag vet allting om dig .
jag kan teckenspråk .
jag känner till proceduren .
jag känner till situationen .
jag lämnade dig ett meddelande .
jag tycker väldigt mycket om Tom .
jag gillar baseboll också .
jag tycker om countrymusik .
jag tycker om ärliga människor .
jag gillar din optimism .
jag ser fram emot det .
jag förlorade medvetandet .
jag tappade bort mina solglasögon .
jag tappade tidsuppfattningen .
jag tycker jättemycket om mitt jobb .
jag gjorde några ändringar .
jag har sociologi som huvudämne .
jag menade tvärtom .
jag träffade Mary i går .
jag missade mötet .
jag måste börja gå hemåt .
jag måste säga någonting .
jag behöver ett större rum .
jag behöver en ny cykel .
jag behöver ett svar nu .
jag behöver lite pengar nu .
jag behöver vägledning .
jag behöver den där medicinen .
jag behöver det där imorgon .
jag måste byta om nu .
jag måste se den nu .
jag måste göra anteckningar .
du måste höra på .
jag behöver era åsikter .
jag behöver dina åsikter .
jag svek dig aldrig .
jag gav aldrig upp hoppet .
jag tyckte aldrig om att gå i skola .
det märkte jag aldrig .
jag litade aldrig på dem .
jag tycker inte om dig längre .
jag beställde pommes frites också .
jag tryckte av .
det där behövde jag verkligen .
jag behövde verkligen det där .
jag behövde verkligen det här .
det här behövde jag verkligen .
jag känner igen den där killen .
jag sade att jag inte var upptagen .
jag såg ett tillfälle .
jag såg en möjlighet .
jag såg dig flina .
jag skickade ett mejl till dig .
jag tvivlar starkt på det .
jag borde antagligen gå .
jag löste mysteriet .
jag löste problemet .
jag fattar fortfarande inte .
jag kommer ännu ihåg Tom .
jag tar danslektioner .
jag tror att Tom ljuger .
jag tror att han var arg .
jag tror att vi borde gå .
jag tror att vi borde åka .
jag tror att du är färdig .
jag tror att ni är färdiga .
jag trodde att jag kände dig .
jag trodde att du åkt .
jag berättade sanningen för Tom .
jag sa det till dig igår .
jag förstår helt och hållet .
jag vill ha någonting nytt .
jag vill dricka mjölk .
jag vill gå till stan .
jag ville träffa dig .
jag ville rädda dig .
jag ville solbada .
jag ville varna Tom .
jag har alltid varit en ensamvarg .
jag höll på att bli sömnig .
jag tittade på henne .
jag var på väg hem .
jag spelade tennis .
jag var väldigt nöjd .
jag hade verkligen otur .
jag var mycket imponerad .
jag blev väldigt överraskad .
jag tvättade fönstren .
jag gick på medicinska fakulteten .
jag önskar dig lycka till .
jag önskar er lycka till .
jag går inte till skolan .
jag tänker inte gå till skolan .
jag skulle inte rekommendera det .
jag skulle inte rekommendera den .
det skulle jag inte gilla .
jag skulle inte gilla det .
jag vore väldigt tacksam .
jag vore mycket tacksam .
det är bäst att jag stannar hemma .
jag skulle vilja vara ensam .
jag skulle vilja följa med dig .
jag skulle vilja se det .
jag skulle vilja stå upp .
jag skulle vilja pröva det här .
jag skulle inte rekommendera det .
jag gör det helst inte .
jag skulle hellre slippa göra det .
jag väntar hellre här .
jag kommer alltid att behöva dig .
jag kommer alltid att behöva er .
jag är tillbaka till dess .
jag kommer att vara tillbaka till dess .
jag kommer tillbaka i tid .
jag är på mitt kontor .
jag kommer att vara på mitt kontor .
jag ringer min man .
jag kommer att drömma om dig .
jag kör dig dit .
jag kör dit dig .
jag kör er dit .
jag kör dit er .
jag skjutsar dig dit .
jag skjutsar dit dig .
jag skjutsar er dit .
jag skjutsar dit er .
jag tar reda på det själv .
jag hämtar Tom åt dig .
jag skall gå till stranden .
jag ska gå till stranden .
jag ska till stranden .
jag tar hand om det här .
jag tar hand om den här .
jag hör av mig .
jag håller dig informerad .
jag håller dig à jour .
jag ska ringa några samtal .
jag kommer att sakna det här stället .
vi ses på jobbet .
vi ses på arbetet .
jag skickar en räkning .
jag skickar en faktura .
jag stannar i bilen .
jag tar en taxi hem .
jag tar chansen .
jag tar tillfället .
jag berättar för de andra .
jag ska berätta för de andra .
jag ska försöka att hitta Tom .
jag kommer att vänta i bilen .
jag väntar på dig .
jag väntar på er .
jag är Marys pojkvän .
jag ringer polisen .
jag väntar ett samtal .
jag är extremt hungrig .
jag känner mig illamående .
jag är färdig med den .
jag är färdig med det .
jag tänker ge den till Tom .
jag tänker ge det till Tom .
jag ger den till Tom .
jag ger det till Tom .
jag är glad att jag hittade dig .
jag är glad att jag hittade er .
jag är glad att det är gjort .
jag är glad att det är över .
jag är glad att du lade märke till det .
jag är glad att du uppmärksammade det .
jag är glad att du märkte det .
jag är glad att du berättade för mig .
jag är glad att ni berättade för mig .
jag är glad att du är här .
jag ska till gymmet .
jag går till gymmet .
jag åker till gymmet .
jag är så gott som aldrig hemma .
jag är nästan aldrig hemma .
jag är här varje kväll .
jag är här för att hjälpa dig .
jag är här för att hjälpa er .
jag är väldigt motiverad .
jag är ytterst motiverad .
jag är kär i dig .
jag ligger i luftvapnet .
jag skämtar med dig bara .
jag skämtar med er bara .
jag driver bara med dig .
jag driver bara med er .
jag driver med dig bara .
jag skojar bara med dig .
jag skojar bara med er .
jag söker arbete .
jag har tur som är här .
jag ska flytta tillbaka hem .
jag är inte hungrig längre .
jag är inte ett dugg trött .
jag undviker inte dig .
jag undviker inte er .
jag är inte upptagen längre .
jag följer inte med .
jag förnekar inte det .
jag kommer inte att dö .
jag ska inte dö .
jag ignorerar dig inte .
jag tänker inte gifta mig med dig .
jag är inte redo att dö .
jag är inte beredd att dö .
jag hindrar dig inte .
jag hindrar er inte .
jag tänker inte hindra er .
jag är inte så synisk .
jag är inte så orolig .
jag har inte på mig det där .
jag har inte på mig den där .
jag tänker inte ha på mig den där .
jag tänker inte ha på mig det där .
jag tänker inte ha på mig det här .
jag tänker inte ha på mig den här .
jag har inte på mig det här .
jag är inte din bror .
jag är inte er bror .
jag är på fel buss .
jag sitter på fel buss .
jag är öppen för vad som helst .
jag är stolt över er alla .
jag är stolt över er allihop .
jag är redo om du är det .
jag är redo om ni är det .
jag är redo att gå vidare .
jag är redo att fortsätta .
jag är ledsen för det här .
jag är tre timmar bort .
jag delar gärna .
jag är villig att dela .
jag är beredd att dela .
jag kan gå med på att dela .
jag arbetar här nu .
jag skriver ett brev .
jag är yngre än Tom .
jag är din nya partner .
jag har varit överallt .
jag har precis ätit middag .
jag har nyss ätit middag .
det har jag aldrig gjort .
jag har aldrig behövt den .
jag har aldrig behövt det .
Imponerande , eller hur ?
är det någon där ?
är det någon där ute ?
är det så illa ?
är det min tur att betala ?
finns det hiss ?
är inte det där Toms hatt ?
är inte det sanningen ?
allt ordnade sig .
det kan inte vara så illa .
det kan vara ett vapen .
den måste avlägsnas .
det är inte Toms fel .
det är inte alltid lätt .
det liknar en anka .
det betyder mycket för mig .
det måste vara ett misstag .
det hela var en stor lögn .
det var ett insidejobb .
det var ett internt jobb .
det var hemskt roligt .
det var inte med vilje .
det hade varit roligt .
det skulle ha varit roligt .
det är 99,9 procent effektivt .
det är nittionio komma nio procent effektivt .
Tom står näst på tur .
det är ett svårt jobb .
det är rena grekiskan för mig .
det är rena rama grekiskan .
för mig är det rena grekiskan .
allt är Toms fel .
det är ett extremfall .
det är kul att titta på tv .
det är skönt att vara tillbaka .
den är gjord av läder .
den är gjord av skinn .
det är skönt att vara hemma .
det angår inte mig .
det står på schemat .
det är ganska spännande .
det är tyst , du vet .
det är middagsdags .
den är värd en förmögenhet .
blunda bara .
ge mig pistolen bara .
hur rik är Tom egentligen ?
sänk rösten .
var snäll och släpp mig .
släpp handtaget .
får jag se den där listan .
låt mig ta en titt .
gör lite nytta .
många av oss är upprörda .
Mary kom självmant .
Mary kom själv .
får jag ställa en fråga ?
får jag låna en linjal ?
kanske jag kan hjälpa till .
kanske jag kan hjälpa dig .
kanske jag kan visa dig .
kanske jag borde göra det .
han kanske inte är ung .
alla män är likadana .
det gör jätteont i min arm .
min chef är väldigt trevlig .
jag fryser om öronen .
min far är frisk .
mina händer skakar .
min mamma är hemma .
mina föräldrar är där .
mina söner är soldater .
inga nyheter är goda nyheter .
ingen har något problem .
ingen har röstat ännu .
ingen är så lycklig .
det var ingen som lyssnade .
ingen hörde på .
ingen kommer att få reda på det .
ingen går in dit .
det är ingen som lyssnar på mig .
ingen behöver tala .
inget av det där spelar någon roll .
ingenting av det här är verkligt .
inget av det här är äkta .
inget av detta är verkligt .
ingenting av det här är sant .
inget av det här är sant .
inget av detta spelar någon roll .
ingenting jag gjorde hjälpte .
inget jag gjorde hjälpte .
ingenting kan gå fel .
inget kan gå fel .
inget här är mitt .
ingenting här är mitt .
ge mig nycklarna nu .
ge mig listan nu .
låt oss komma igång .
okej allesamman , hör på nu .
okej allihopa , hör på .
en av dem ljuger .
en av dem var min .
ett av dem var mitt .
spela den sången igen .
var snäll och ta med en sallad .
kaniner tycker om morötter .
kaniner gillar morötter .
Room service , tack .
Rumsservice , tack .
hon tillät mig gå .
hon brast i gråt .
hon har tio barn .
han är min vän .
hon är min flickvän .
hon vill döda mig .
hon blev påkörd av en bil .
hon kommer förmodligen .
borde jag klippa mig ?
borde jag klippa håret ?
ska jag öppna den nu ?
Storleken har ingen betydelse .
så vad betyder det ?
ta en titt på de här .
ta en titt där inne .
säg åt Mary att jag älskar henne .
säg till Tom att det är brådskande .
säg åt Tom att skriva till mig .
berätta för mig hur man gör .
berätta för mig hur jag ska göra .
berätta vad du såg .
det var inte överenskommelsen .
det där var inte överenskommelsen .
det var inte planen .
det där är Toms teckning .
det är väldigt personligt .
det är där jag kommer att vara .
dörren är öppen nu .
hela gänget är här .
garaget var tomt .
hästen hoppar .
huset brinner .
huset står i brand .
Mjölken kokade över .
Apan kom ner .
den gamle mannen satte sig ner .
telefonen ringer .
telefonen ringde igen .
Talaren är ung .
texten är för lång .
vinden avtog .
det finns villkor .
det finns en fågel här .
det finns ingen lösning .
det finns en krona här .
det är en krona här .
det står ett glas här .
det finns ett glas här .
de här är de enda jag har .
de närmar sig .
de är vegetarianer .
det sade de inte .
det sa de inte .
de bor på nedre våningen .
de började dansa .
de gick ut .
de sade åt oss att vänta .
de var sårbara .
de ville inte lyssna .
de är alla barfota .
de är barfota allihop .
de är barfota allesammans .
de är där inne allihop .
de är där inne allesammans .
de är likadana allihop .
de är likadana allesammans .
de är svåra att hitta .
de är på mitt kontor .
de är inte hemma än .
det är inte mina regler .
det här måste upphöra .
det här måste få ett slut .
det här är Toms skola .
detta är Toms skola .
det här är en bra början .
det här är en jättebra idé .
det här är en trollstav .
det här är en säker plats .
det här är en liten bok .
det här börjar bli svårt .
detta är vårt beslut .
detta är inte acceptabelt .
det här är mycket allvarligt .
det här handlar inte om dig .
detta handlar inte om dig .
det här handlar inte om er .
detta handlar inte om er .
den här måste vara till dig .
den här pennan är bäst .
den här mattan är handgjord .
det är våra order .
Tom kan inte vara allvarlig .
Tom kan inte vara seriös .
Tom kollade datumet .
Tom kollade tiden .
Tom kunde inte hacka den .
Tom kunde inte hacka sig in i den .
Tom kunde inte hjälpa oss .
Tom hann inte med .
Tom klarade sig inte .
Tom kunde inte komma .
Tom kräver uppmärksamhet .
Tom har behov av uppmärksamhet .
Tom gjorde ett halv @-@ färdigt jobb .
Tom dödade inte Mary .
Tom kände inte Mary .
Tom såg inte upptagen ut .
Tom äter inte kött .
Tom får inte betalt .
Tom hatar dig inte .
Tom hatar er inte .
Tom hatar inte dig .
Tom hatar inte er .
Tom drack i tystnad .
Tom har hjälpt till mycket .
Tom har varit till stor hjälp .
Tom har många talanger .
Tom har dålig hygien .
Tom har tre farbröder .
Tom har tre morbröder .
Tom har inte mått bra .
Tom har inte ringt mig .
Tom är miljardär .
Tom är lite udda .
Tom är lite konstig .
Tom är brandman .
Tom är en bra vän .
Tom är en bra person .
Tom är neurolog .
Tom är nervspecialist .
Tom är redan där .
Tom är annorlunda nu .
Tom sitter i fängelse nu .
Tom är i duschen .
Tom är precis som du .
Tom är lång och smal .
Tom tittar på den .
Tom tittar på mig .
Tom ser trött ut .
Tom kommer aldrig i tid .
Tom är väldigt charmig .
Tom är inte en trevlig kille .
Tom är inte en sympatisk kille .
Tom är inte en schyst kille .
Tom är inte någon schyst kille .
Tom är ingen främling .
Tom är inte stor nog .
Tom är inte tillräckligt stor .
Tom ligger inte ned .
Tom säger inte varför .
Tom är inte så säker .
Tom är inte så galen .
Tom försvann just .
Tom försvann bara .
Tom försvann precis .
Tom gick just in .
Tom gick bara in .
Tom visste att jag hade rätt .
Tom slog ner honom .
Tom vet att han har rätt .
Tom vet att vi är här .
Tom lät Mary gå hem .
Tom gillar reality @-@ tv .
Tom tycker om reality @-@ tv .
Tom ser skräckslagen ut .
Tom ser frustrerad ut .
Tom ser väldigt glad ut .
Tom gjorde en bra putt .
Tom lovade att hjälpa .
Tom sade att han berättat för dig .
Tom sade att han berättat för er .
Tom säger sig vara hungrig .
Tom halkade och föll .
Tom låter utmattad .
Tom började klättra .
Tom började skratta .
Tom stal dina pengar .
Tom stal era pengar .
Tom simmade i simbassängen .
Tom tror att jag har rätt .
Tom tycker att jag har rätt .
Tom sade att Mary skulle ljuga .
Tom sade att jag skulle göra det .
Tom sade åt mig att köra .
Tom försökte döda mig .
Tom försökte rädda mig .
Tom snavade och föll .
Tom avrättades i elektriska stolen .
Tom gavs en dödande elektrisk stöt .
Tom var inte borta länge .
Tom var inte förvånad .
Tom var inte särskilt upptagen .
Tom gick ut och dansade .
Tom kommer att bli överlycklig .
Tom kommer inte att komma i tid .
Tom gav sig inte .
Tom gav inte vika .
Tom skulle inte ge sig .
Tom skulle inte ge vika .
Tom fötter kändes stelfrusna .
Tom hade ingen känsel i fötterna .
Tom börjar bli frusen .
Tom är min vän med .
Tom är min vän också .
försök att inte vara dum .
försök vara modig , Tom .
försök att komma på det .
försök komma på det .
var han fallskärmsjägare ?
vi visste alla om det .
vi visste alla om den .
vi jobbar alla för hårt .
vi tar alltid bussen .
vi äter middag .
vi är inte amerikaner .
vi kan alla gå hem .
vi kan beställa pizza .
vi kan ännu göra det .
vi kan prata om det .
vi kan behöva din hjälp .
kan vi lösa det här ?
vi kan inte gå in dit .
vi pratade om det .
vi har ett trevligt hus .
vi har saker att göra .
vi måste göra bättre ifrån oss .
vi måste lämna dig .
vi måste få ett slut på det här .
vi måste berätta det för dem .
vi måste vänta här .
vi har två barn .
vi har jobb åt Tom .
vi hoppas att det här är sant .
vi hoppas att det här stämmer .
vi matade just babyn .
vi matade just barnet .
vi kysstes .
vi visste allt om det .
vi visste allt om den .
vi behöver ett säkerhetsnät .
vi behöver hjälp här inne .
vi måste vila oss snart .
vi måste prata mera .
vi måste vänta här .
vi borde sätta upp en fälla .
vi reste tillsammans .
vi tittar på tv tillsammans .
vi gick till stranden .
vi var alla så trötta .
vi var nästan där .
du tänkte försöka .
vi höll på att äta lunch .
vi skulle just gå .
vi lekte bara .
vi hade delvis rätt .
vi var ganska högljudda .
vi förde ganska mycket oljud .
vi var väldigt nära varandra .
vi stannade uppe hela natten .
vi jobbade sent .
vi skickar det till dig .
vi träffar Tom senare .
vi möter dig där .
vi möter er där .
vi hämtar dig där .
vi hämtar er där .
vi är extremt upptagna .
vi är vänner , eller hur ?
vi är i en konjunktursvacka .
vi är i en recession .
vi är i en lågkonjunktur .
vi är inte så nära .
vi är redo för detta .
vi är oentusiastiska .
vi har listat ut det .
vilken kreativ idé !
vilken trevlig överraskning !
vilken märklig kvinna !
vilken underlig kvinna !
vilken fantastisk idé !
vad har du för alternativ ?
vad säger de ?
vad lagar du ?
vad ska du ta ?
vad tvättar du ?
vad har du på dig ?
vad har du på dig för kläder ?
vad skriver du ?
vad för dig hit ?
vad kan du ge mig ?
vad kan du ge oss ?
vad kan du berätta för oss ?
vad kan du tala om för oss ?
vilken färg var de ?
vad kunde det betyda ?
vad snubblade jag på ?
vad kallade Tom mig för ?
vad gjorde Tom här ?
vad gjorde Tom sedan ?
vad föreslog Tom ?
vad sade han till dig ?
vad sade han till er ?
vad berättade han för dig ?
vad berättade han för er ?
vad betydde allt det där ?
vad gjorde vi fel ?
vad frågade du av Tom ?
vad kallade du mig ?
vad kallade ni mig ?
vad gjorde du sedan ?
vad gav du upp ?
vad har du grävt fram ?
vad har vi här ?
vad vill vi här ?
vad känner du nu ?
vad minns du ?
vad minns ni ?
vad bevisar det ?
vad mer kan jag förlora ?
vad mer kan du göra ?
vad mer kan ni göra ?
vad annat har vi ?
vad annat behöver vi ?
vad annat ser du ?
exakt vad är det där ?
vad är det som pågår här inne ?
vilken årskurs är Tom i ?
vad bör jag göra nu ?
vad var Toms brott ?
vad ska jag säga till Tom ?
vad är det du räknar ?
vad räknar du ?
vad är det ni räknar ?
vad räknar ni ?
vad tittar du på ?
vad tittar ni på ?
vad är Toms problem ?
vad är det i korgen ?
vad finns i garderoben ?
vad är det i kaffet ?
vad står på dagordningen ?
vad har du på tallriken ?
vad är planen , Tom ?
vad är deras syfte ?
vad är syftet med dem ?
vad är ditt smeknamn ?
vad är din lösning ?
vad är er lösning ?
när frågade du Tom ?
när kom du in ?
när gjorde du det ?
när gjorde du det här ?
när gav du upp ?
när såg du Tom ?
när talade du om det för mig ?
när behöver de mig ?
när ska Tom vara tillbaka ?
när kommer du tillbaka ?
var är hästarna ?
var är polisen ?
vart är vi på väg ?
vart är du på väg ?
var kan jag hitta Tom ?
var kan jag träffa Tom ?
var köpte Tom den ?
var har du fått det ifrån ?
var satte du den ?
var hittar jag det ?
var är hennes bild ?
var ligger tvättstugan ?
var är tvätten ?
var är din jacka ?
var ligger er skola ?
var är ingången ?
var är tvättrummet ?
var är ditt bagage ?
var är ert baggage ?
var är era bagage ?
vem kan jag sälja den till ?
vem kan utföra det här arbetet ?
vem röstade du på ?
vem tycker inte så ?
vad annat saknar du ?
vem annan är där inne ?
vem mer är därinne ?
vem mer är där inne ?
vem annan var här inne ?
vem sa att jag har en pistol ?
vem satt här ?
vem skrev brevet ?
vem är redo att beställa ?
varför är ni alla här ?
varför gör du det ?
varför är du här nu ?
varför är du hemma nu ?
varför känner du dig kränkt ?
varför sover du ?
varför är du så nervös ?
varför är du så trött ?
varför är de inte tillbaka ?
varför är inte de tillbaka ?
varför är de inte här ?
varför är inte de här ?
varför är du inte där ?
varför är ni inte där ?
varför är inte du där ?
varför är inte ni där ?
varför ringde Tom till dig ?
varför sa Tom det ?
varför sa Tom så ?
varför tog du med den ?
varför köpte du den där ?
varför köpte du det där ?
varför sparkade du Tom ?
varför avskedade du Tom ?
varför lämnade du oss ?
varför valde du Tom ?
varför sköt du mig ?
varför talade du om det för Tom ?
varför har du den där ?
varför har du den här ?
varför behöver du den här ?
varför stannar du här ?
varför vill du ha det där ?
varför gör Tom det där ?
varför svarar du inte ?
varför sover inte Tom ?
varför var inte Tom där ?
igår var det måndag .
igår var det söndag .
du ljuger alltid för mig .
du kan komma in igen .
du kan komma in här .
du kan ordna allt det här .
du kan börja gå hemåt .
du kan hålla min hand .
du kan åka med mig .
du kan sitta ned nu .
du kan sätta dig nu .
ni kan sitta ned nu .
ni kan sätta er ned nu .
du kan stanna här inne .
du kan stanna hos mig .
du kan stanna hos oss .
du kan använda min telefon .
du kan inte ändra på Tom .
ni kan inte ändra på Tom .
man kan inte ändra på Tom .
du kan inte kontrollera mig .
ni kan inte kontrollera mig .
man kan inte kontrollera mig .
du kan inte följa med oss .
du kunde ha sagt nej .
du skulle kunna sagt nej .
du skulle kunna ha sagt nej .
du förstår inte .
ni förstår inte .
du gav mig för mycket .
du gav upp för fort .
du får ta nästa .
du kom undan med det .
du hann hit i tid .
du hann hit i tid .
du har missförstått det hela .
du har ett jättebra jobb .
du måste vara redo .
du måste välja en .
du måste välja ut en .
du måste berätta för Tom .
du måste berätta det för Tom .
du måste lita på mig .
ni måste lita på mig .
du måste prova det här .
du måste försöka , Tom .
du vet att jag kan göra det .
du vet att jag klarar det .
du måste vara så stolt .
du måste göra som jag säger .
ni måste göra som jag säger .
du måste komma hem .
du måste hjälpa Tom .
du behöver det jag har .
du verkar hata Tom .
ni verkar hata Tom .
du är en bra doktor .
du är en bra läkare .
du är duktig på att kyssas .
du är en bra sångare .
du är lite sen .
ni är lite sena .
du är en soldat nu .
du är allt de har .
du är allt som de har .
ni är allt de har .
ni är allt som de har .
ni är alla väldigt lugna .
du är nästa trettio .
ni är nästan trettio .
du är en timme tidig .
ni är en timme tidiga .
du är ohövlig .
du är respektlös .
ni är oansvariga .
du är inte misstänkt .
det är inte du som bestämmer .
du är vårt enda hopp .
du är överkänslig .
ni är överkänsliga .
du har verkligen talang .
ni har verkligen talang .
du är så bra på det .
ni är så bra på det .
du är för lättsinnig .
du är oberäknelig .
ni är oberäkneliga .
du är väldigt flexibel .
du är väldigt vig .
du har gjort rätt .
ni har gjort rätt .
din hund bet mig i handen .
talar jag för snabbt ?
pratar jag för snabbt ?
vad som helst blir bra .
är muffinsen färdiga ?
finns det några bananer ?
är det där mina örhängen ?
är du en riktig läkare ?
njuter du av det här ?
njuter du av detta ?
njuter ni av det här ?
njuter ni av detta ?
är du road av det här ?
är du road av detta ?
är ni roade av det här ?
är ni roade av detta ?
väntar du på Tom ?
stöter du på mig ?
är du hungrig över huvud taget ?
är du fortfarande hemma ?
är ni fortfarande hemma ?
är du fortfarande gift ?
är ni fortfarande gifta ?
är ni två musiker ?
bananer är goda .
kan du stanna en minut ?
kan du inte röra dig fortare ?
katter tycker inte om vatten .
skulle jag kunna få en servett ?
skadades någon ?
köpte ni Tom en hund ?
köpte du en hund till Tom ?
köpte ni en hund till Tom ?
köpte du en ny bil ?
köpte ni en ny bil ?
kom du med tåget ?
åt du frukost ?
åt ni frukost ?
ringde du någonsin Tom ?
fick du checken ?
fick ni checken ?
kände du Tom väl ?
kände ni Tom väl ?
tror du på mig nu ?
tror ni på mig nu ?
blir du någonsin snurrig ?
blir ni någonsin snurriga ?
flyger du ofta ?
flyger ni ofta ?
måste du gå nu ?
måste ni gå nu ?
måste ni åka nu ?
måste du åka nu ?
tycker du om ansjovis ?
gillar du sött te ?
tycker du om den här staden ?
tycker du om att resa ?
menar du det på riktigt ?
Jaså , menar du det ?
talar du japanska ?
älskar du honom fortfarande ?
tycker du att jag är ful ?
tycker ni att jag är ful ?
använder du aftershave ?
använder ni aftershave ?
använder du rakvatten ?
spelar det verkligen någon roll ?
talar hon franska ?
prata inte ens med mig .
tala inte ens med mig .
förvänta dig inte övertid .
glöm inte att använda tandtråd .
glöm inte din väska .
ge inte upp halvvägs .
låt inte Tom se dig .
låt inte Tom se er .
låt inte Tom vissla .
se inte så chockad ut .
Tvinga mig inte att göra detta .
Tvinga mig inte att göra det här .
för inte oväsen här .
öppna inte fönstret .
peka inte på andra .
svara inte på det .
Stirra inte på folk .
Ödsla inte din tid .
Ödsla inte er tid .
slösa inte bort er tid .
Maska inte .
Dubbelklicka på ikonen .
ät vad du vill .
ät vad ni vill .
ät vadhelst du vill .
ät vadhelst ni vill .
Europa är en kontinent .
alla var ängsliga .
allt blev svart .
allting blev svart .
allt förändras .
fyll i den här , tack .
fyll i denna , tack .
Lyckan log mot honom .
det är rea på pälskappor .
ge mig det där kuvertet .
ge mig tre minuter .
ge oss tre minuter .
glad alla hjärtans dag .
har de kommit än ?
har du rökt ?
har du sett Tom än ?
har ni sett Tom än ?
han beundrade min nya bil .
han gör alltid anteckningar .
han frågade mig vem jag var .
han blev polis .
han kom för sent som vanligt .
han gav mig ett exempel .
han har en massa böcker .
han har många böcker .
han har massor av böcker .
han är alltid punktlig .
han är bra på att sjunga .
han är bara en amatör .
han är inte alltid sen .
han är inte snäll mot henne .
han tvättar bilen .
han har på sig glasögon .
han tycker mycket om fotboll .
han gifte sig med en skådespelerska .
han rånade en gammal dam .
han satt och läste en bok .
han vände sig i sängen .
han blev exkommunicerad .
han är en riktig gentleman .
han är modig och ärlig .
han går upp tidigt .
han stiger upp tidigt .
han kliver upp tidigt .
han är inte alltid glad .
han berättelse låter sann .
hans historia låter sann .
hur upptagen kan Tom vara ?
hur vet du det ?
hur vet ni det ?
hur gjorde du det ?
hur gjorde ni det ?
hur visste Tom det ?
hur träffade Tom Mary ?
hur kom du dit ?
hur tog du dig dit ?
hur fick du tag på dem där ?
hur mjölkar man en ko ?
hur länge var Tom här ?
vad kostar det ?
hur gammal är din morbror ?
jag skördar vete .
jag uppskattar hjälpen .
jag antog att det var gratis .
jag antog att den var gratis .
jag blev Toms vän .
jag lånade Toms cykel .
jag köpte den i går .
jag kom hem sent .
jag kom hit i går .
jag kan inte äta choklad .
jag hittar inte mina skor .
jag hör ingenting .
jag får inte upp den här burken .
jag kommer hit varje dag .
jag skulle kunna få henne att prata .
jag kunde inte ljuga för dig .
jag kunde inte ljuga för er .
jag fick inte hyra en bil .
jag bad inte om detta .
jag bad inte om det här .
jag förstod inte hans skämt .
jag gick inte till skolan .
jag flyttade inte på någonting .
jag sade inte att jag höll med .
jag sa inget .
jag sa ingenting .
jag ogillar att vara ensam .
jag får inte så mycket post .
jag vet inte vem jag är .
jag gillar ingenting .
jag behöver ingen hjälp .
jag pratar inte svenska .
jag talar inte svenska .
jag vill inte tillbaka .
jag vill inte ha något vin .
jag vill inte ha dig här .
jag vill inte ha er här .
jag konstaterade en sak .
jag fick reda på någonting .
jag kom underfund med någonting .
jag får åksjuka .
jag åker dit varje år .
jag blev blöt ända in på skinnet .
jag var tvungen att göra någonting .
jag är kär i dig .
jag svärmar för dig .
jag har några funderingar .
jag har några tankar .
jag har några idéer .
jag har en halvbror .
jag har en förklaring .
jag har ett till alternativ .
jag har ett alternativ till .
jag har ett annat alternativ .
jag har tappat bort min plånbok .
jag har inga pengar på mig .
jag har tre barn .
jag måste gå och sova .
jag fick precis ditt mejl .
jag fick precis ditt mail .
jag stötte precis min tå .
jag stötte precis tån .
jag visste att jag inte var galen .
jag kände alla där .
jag visste vad du menade .
jag visste vad ni menade .
jag känner Tom personligen .
jag vet hur gammal Tom är .
jag vet hur detta fungerar .
jag vet hur det här funkar .
jag gillar hur Tom tänker .
jag tycker om hur Tom tänker .
jag tycker om att spela tennis .
jag gillar att vara förberedd .
jag tycker om att spela tennis .
jag älskar att spela Chopin .
jag älskar att prata med dig .
jag älskar att prata med er .
jag stavade fel på ordet .
jag måste bege mig nu .
jag måste ge mig av nu .
jag måste göra min läxa .
jag måste ha drömt det .
jag behöver den i morgon .
jag behöver den till i morgon .
jag måste bädda min säng .
jag behöver att du går hem .
jag fick aldrig veta varför .
jag gick aldrig och lade mig .
jag övade varje dag .
jag satte Tom på listan .
jag kommer ihåg den kvällen .
jag säger det hela tiden .
jag nyser hela tiden .
jag gillar det fortfarande inte .
jag tycker fortfarande inte om det .
jag berättar allt för Tom .
jag tror att Mary tycker om mig .
jag tror att Mary gillar mig .
jag tror inte att han kommer .
jag tror att det är en bluff .
jag trodde att jag hörde dig .
jag trodde att jag var ensam .
jag trodde att jag var lyckligt .
jag tyckte att jag var lycklig .
jag tyckte att det var gott .
jag tyckte att det var bra .
jag trodde att du skulle hålla med .
jag brukade spela tennis .
jag vill att Tom går hem .
jag vill att Tom åker hem .
jag vill ha något annat .
jag vill tro dig .
jag vill tro er .
jag vill tillbaka nu .
jag vill följa med dig .
jag hade inte bråttom .
jag var inte alltför trött .
jag kommer att behöva din hjälp .
jag ska skriva om det .
jag tänker skriva om det .
jag önskar att jag hade ringt Tom .
jag önskar att du skulle ringa Tom .
jag kommer inte att låta det hända .
jag kommer inte att göra någon polisanmälan .
jag kommer inte stanna hos dig .
jag undrar varför Tom stack .
jag undrar varför Tom drog .
jag undrar varför Tom åkte .
jag undrar varför Tom gick .
jag arbetar på ambassaden .
jag skulle ha skickat rosor .
jag skulle inte ljuga för dig .
jag skulle inte ljuga för er .
jag skulle inte ta i den där .
jag skulle gå med på att betala .
jag skulle vara villig att betala .
jag skulle vara beredd att betala .
det är bäst att jag rör på mig .
jag skulle göra likadant .
jag skulle göra samma sak .
jag skulle dubbelkolla det .
jag skulle dubbelkontrollera det .
jag skulle känna likadant .
jag skulle vilja samarbeta .
jag skulle vilja gå in .
det skulle jag vilja höra .
jag skulle aldrig drömma om det .
jag skulle hellre vara och fiska .
jag bor hellre ensam .
jag skulle säga att du förtjänade det .
jag skulle säga att du gjorde dig förtjänt av det .
jag skulle fortfarande vilja försöka .
jag skulle fortfarande vilja pröva .
jag ringer honom ikväll .
jag ringer honom i kväll .
jag hämtar den åt dig .
jag hämtar det åt dig .
jag kommer till saken .
jag går om du insisterar .
jag kommer snart träffa honom
jag går och tvättar händerna .
jag ska ringa några samtal .
jag kommer aldrig att förstå .
jag ska tänka på det .
jag försöker att få tag i Tom .
jag försöker att nå Tom .
jag är lite uppskakad .
jag är rädd för höjder .
jag är inte rädd för någonting .
jag är rädd för spindlar .
jag är rädd för att gå hem .
jag är rädd för att åka hem .
jag är nästan säker på det .
jag är vid den norra porten .
jag är vid den norra grinden .
jag är trött på Boston .
jag ringer Tom igen .
jag är bekväm med det
jag gör mina läxor .
jag är glad att jag fångade dig .
jag är glad att jag var i närheten .
jag är glad att vi hittade dig .
jag är glad att vi hittade er .
jag är glad att du gillar Tom .
det gläder mig att du tycker om Tom .
det gläder mig att du kommer ihåg .
det gläder mig att du minns .
det gläder mig att ni minns .
det gläder mig att ni kommer ihåg .
jag är glad att du är tidig .
jag är glad att ni är tidiga .
jag går tillbaka till sängen .
jag går tillbaka till sängs .
jag är här för att be om ursäkt .
jag är bara ärlig .
jag känner mig bara nere .
jag är ledig från arbetet i morgon .
jag är säker på att det inte är någonting .
jag har varit sämre .
jag har varit upptagen .
jag har varit ganska upptagen .
jag har varit där mycket .
jag har lånat ett bord .
jag har massor att göra .
jag har massvis med saker att göra .
jag har några kakor .
jag har precis kommit hem .
jag har sett det här förut .
jag har sett detta förut .
jag har slutat räkna .
jag har slutat att räkna .
är det din egen idé ?
stämmer inte det , Tom ?
eller hur , Tom ?
är inte det misstänksamt ?
är inte svaret lätt ?
det regnar kraftigt .
det gjorde ingen skillnad .
det påminde mig om dig .
det påminde mig om er .
det är helt klart lämpligt .
det var förståeligt .
det var begripligt .
det var väldigt svårt .
det var inte mitt beslut .
det var inte sensationellt .
det var inte uppseendeväckande .
det var inte fantastiskt .
det är måndag , du vet .
den är kvart i två .
det är fullständigt fel .
det är en omöjlighet .
det har varit intressant .
det är för barnen .
det är till barnen .
det är mitt jobb , du vet .
det är inte akut .
det är ingenting personligt .
det är troligen hemsökt .
det är troligtvis hemsökt .
det är antagligen hemsökt .
det spökar troligtvis där .
det är verkligen vackert .
den är verkligen vacker .
det är för överväldigande .
det är väldigt intressant .
det är ditt val , Tom .
Jesus var snickare .
ett ögonblick .
andas bara som vanligt .
gå inte ut bara .
ge oss en minut bara .
håll Tom utanför detta .
håll Tom utanför det här .
släpp in lite frisk luft .
låt mig fråga en fråga .
låt mig ställa en fråga .
låt mig ringa min advokat .
låt mig ta hand om Tom , okej ?
låt mig tänka en minut .
låt mig fundera en minut .
kärlek är för tonåringar .
Markera rätt svar .
Mary är en gold @-@ digger .
Maj kommer efter april .
min katt dog i går .
min mor älskar musik .
mitt rum är mycket litet .
ingen skulle skada Tom .
ingen skulle ha brytt sig .
ingen här äter kött .
ingen anmäler sig frivilligt .
ingen ställer upp frivilligt .
inte alla fåglar kan flyga .
det är inte alla fåglar som kan flyga .
ingenting hände här .
varför är du här ?
Optimister lever längre .
var snäll och dela ut korten .
var snäll och stryk skjortan .
Ställ undan cykeln .
var inte orolig .
hon skyndade ner för trapporna .
hon följde honom hem .
hon har en fin docka .
hon strök hans skjortor .
hon är en god simmare .
hon är lika lång som du .
hon måste hjälpa honom .
hon tog sitt liv .
borde inte du gå hem ?
borde inte ni gå hem ?
borde inte du åka hem ?
borde inte ni åka hem ?
så vart ska ni ?
så vart ska du ?
så vart ska ni åka ?
så vart ska du åka ?
så vart ska du gå ?
så vart ska ni gå ?
någon tappade sin plånbok .
någon tappade en plånbok .
sluta vara så nyfiken .
sluta jämra dig !
studera de här meningarna .
ta väl hand om Tom .
berätta för mig vad Tom sa .
säg mig vad jag ska tänka .
tack för allt .
tack för ditt svar .
tack för ert svar .
den där mannen är en soldat .
det är rätt åt honom .
rätt åt dig !
det var Toms mamma .
det där var Toms mamma .
det var nära ögat .
det kommer att göra mig lycklig .
det är bara en ursäkt .
det är en del av mitt arbete .
det är förmodligen säkrare .
det är deras angelägenhet .
spädbarnet log mot mig .
isen är väldigt tjock .
Pajen smakade utsökt .
dammen har torkat ut .
soldaterna är döda .
staden var öde .
staden låg öde .
vinden blåste hela dagen .
det blåste hela dagen .
Kvinnorna arbetar .
det är ett par här .
det finns ett par här .
de kunde inte hjälpa oss .
de började skjuta .
de pratade hela natten .
de kommer inte att komma i tid .
de är alla olika .
båda skrattar .
bägge skrattar .
de är tungt beväpnade .
de är inte fångar .
detta är en katastrof .
det här är en snuskig film .
det här är också ett äpple .
detta är också ett äpple .
det här är ett gammalt brev .
detta är ett gammalt brev .
det här är en besvikelse .
det här är inte något misstag .
detta är inte något misstag .
detta är inget misstag .
det här vinet smakar gott .
det här vinet är gott .
det här kommer inte att göra ont alls .
det oroar mig mycket .
Tom bad mig om hjälp .
Tom åt en snabb lunch .
Tom åt en snabblunch .
Tom blev väldigt upprörd .
Tom har inte råd med båda .
Tom har inte råd med bägge .
Tom kan inte ersättas .
Tom kan inte hantera det här .
Tom kan inte stå still .
Tom sprang efter Mary .
Tom skulle kunna vara var som helst .
Tom kunde knappt gå .
Tom stod inte ut med det .
Tom gjorde det , eller hur ?
Tom såg sig inte om .
Tom såg inte tillbaka .
Tom tänkte inte tillbaka .
Tom drog sig inte ur .
Tom backade inte ut .
Tom tycker inte om öl .
Tom bor inte här .
Tom ser inte upptagen ut .
Tom verkar inte upptagen .
Tom kom i vägen för Mary .
Tom hoppade av sin häst .
Tom växte upp på en bondgård .
Tom har en bokning .
Tom har gjort sitt bästa .
Tom lade på telefonen .
Tom la på telefonen .
Tom är Marys skyddsling .
Tom är Marys protegé .
Tom är bilförsäljare .
Tom är en desertör .
Tom är en värnpliktsvägrare .
Tom är en helbrägdagörare .
Tom är en bra make .
Tom är en hemmaman .
Tom är lite galen .
Tom är en urusel dansare .
Tom är på flygplatsen .
Tom är upptagen , eller hur ?
Tom är inte Marys typ .
Tom är inte en bra kock .
Tom är inte heller upptagen .
Tom är inte upptagen heller .
Tom samarbetar inte .
Tom hjälper inte till något .
Tom är inte riktigt säker .
Tom är inte så stark .
Tom är inget ljushuvud .
Tom är inget större ljus .
Tom dödade spindeln .
Tom vet att jag väntar .
Tom kan lite franska .
Tom vet att det är sant .
Tom vet att du är här .
Tom vet att ni är här .
Tom lämnade vattnet på .
Tom ser orolig ut nu .
Tom sänkte rösten .
Tom gjorde många ändringar .
Toms huvudämne var franska .
Tom måste ha haft en nyckel .
Tom behöver vinna tid .
Tom har ofta på sig en hatt .
Tom lade ned boken .
Tom la ner boken .
Tom sprang med full fart .
Tom skakade Marys hand .
Tom tog Mary i hand .
Tom tycker att det är roligt .
Tom tycker att det är kul .
Tom tycker att det är jättebra .
Tom tog Marys ställe .
Tom tog Marys plats .
Tom tog alla mina pengar .
Tom stängde av tv:n .
Tom ville ha mer utrymme .
Tom kommer inte att förlåta dig .
Tom kommer inte att förlåta er .
Tom kommer inte att låta dig betala .
Toms väskor är packade .
Tom är inte alls säker .
Tom är väldigt , väldigt bra .
Tom har fel , vet du .
vänta . skjut inte än .
vi bakar kakor .
vi har inga hemligheter .
vi hör ingenting .
vi hör inget alls .
vi hör ingenting alls .
vi har tre minuter .
vi lyssnar med öronen .
vi behöver bara en minut .
vi visste att Tom skulle vinna .
vi byggde ett sandslott .
vi gjorde ett sandslott .
vi behöver några minuter .
vi behövde information .
vi gick till museet .
vi kommer att behöva deras hjälp .
vi ligger lite efter .
vi är nästan färdiga .
vi är försenade .
vi ligger efter .
vi släpar efter .
vi ligger efter i tid .
vi diskuterar det .
vi är i behov av hjälp .
vi är aldrig nöjda .
vi är inte ansvariga .
vi måste varna Tom .
vi har fått in ett klagomål .
vi fick den analyserad .
vi fick det analyserat .
vi har träffats några gånger .
vi har aldrig behövt det .
vi har aldrig behövt den .
vi har slut på kol .
lyssnade inte du ?
lyssnade inte ni ?
vilken spännande match !
vad är de gjorda av ?
vad anspelar du på ?
vad kan jag göra för dig ?
vad kan jag göra för er ?
vad har du gjort idag ?
vad sa du till Tom ?
vad sa ni till Tom ?
vad berättade du för Tom ?
vad berättade ni för Tom ?
vad mer åt Tom ?
vad mer sa Tom ?
vad mer behöver du ?
vad hände i natt ?
vad händer i morgon ?
vad har du inte gjort ?
vad är Tom rädd för ?
vad är det som pågår här ?
vilket skepp var du på ?
ombord på vilket skepp var du ?
vad gör vi här ?
vad gör Tom här ?
varför gömmer sig Tom ?
vad är det Tom gömmer sig för ?
vad heter hon nu igen ?
vad finns det i den här byrålådan ?
vad finns det i den här lådan ?
vad är det som tar så lång tid ?
vad är det som tar en sådan tid ?
var har du fått det där ärret ifrån ?
var kommer det där ärret ifrån ?
var befinner de sig ?
vad är det för fel på dig ?
när sa Tom det ?
när fick du reda på det ?
när fick du den här ?
när fick ni den här ?
när sa du det ?
när sa ni det ?
när sa du det där ?
när sa ni det där ?
när behöver Tom den ?
när ska uppsatsen lämnas in ?
när är din födelsedag ?
när blir det klart ?
var växte du upp ?
var växte ni upp ?
var bor du nu ?
var bor ni nu ?
var är hissen ?
var är ingången ?
var är skeppet nu ?
var är era bagage ?
var ska jag lägga den ?
var är tidningen ?
var ligger tidningen ?
var är din bil , Tom ?
var är er bil , Tom ?
var är din son , Tom ?
vem talar jag med ?
Vilka är Toms vänner ?
Vilka pratade ni med ?
vem pratade ni med ?
vem pratade du med ?
Vilka pratade du med ?
vem har inte varit där ?
vem uppfann dubbelslipade glasögon ?
vem sålde dig den här bilen ?
vem sålde den här bilen till dig ?
vem skrev det här brevet ?
vem skulle vilja döda mig ?
Vilka gifter sig ?
vems sida är du på ?
på vems sida är du ?
vems sida är ni på ?
vem står näst på tur ?
varför frågar du mig ?
varför sover inte du ?
varför sover inte ni ?
varför sover du inte ?
varför sover ni inte ?
varför kan du inte hjälpa mig ?
varför kan ni inte hjälpa mig ?
varför hatar Tom dig ?
varför hatar Tom er ?
jag kan väl skjutsa dig ?
varför skjutsar inte jag dig ?
varför är Tom här idag ?
varför är tåget sent ?
varför är inte Tom hemma ?
varför sitter inte Tom i fängelse ?
varför sitter inte Tom i häkte ?
varför ler inte Tom ?
varför berättar du inte för oss ?
varför berättar ni inte för oss ?
varför skulle Tom hjälpa oss ?
stannar du hemma ?
ska du resa ensam ?
skulle inte det vara trevligt ?
yoga kommer från Indien .
ni ser alla så glada ut .
ni ser alla så lyckliga ut .
bara du kan göra detta .
mig lurar du inte !
mig lurar ni inte !
man kan inte köpa respekt .
du kan inte köpa respekt .
du kan inte ersätta Tom .
du måste inte äta .
du har många vänner .
du måste gå nu .
du ser så vacker ut .
du måste gå till skolan .
du borde lita på mig .
du verkade lycklig här .
du verkade glad här .
du var inte borta länge .
ni var inte borta länge .
du var inte här då .
ni var inte här då .
du var inte särskilt trevlig .
ni var inte särskilt trevliga .
du skulle ha gillat det .
ni skulle ha gillat det .
du skulle ha tyckte om det .
ni skulle ha tyckt om det .
du skulle inte njuta av det .
du skulle inte tycka om det .
ni skulle inte tycka om det .
ni skulle inte njuta av det .
du skulle inte finna nöje i det .
ni skulle inte finna nöje i det .
du skulle inte tycka om Tom .
ni skulle inte tycka om Tom .
du skulle inte gilla Tom .
ni skulle inte gilla Tom .
du kommer inte att ha något val .
det kommer att missa frukosten .
du är Toms favorit .
du är alltid försiktig .
ni är alltid försiktiga .
du är alltid noggrann .
ni är alltid noggranna .
du beter dig barnsligt .
du hör saker .
nu mumlar du igen .
ni är inte så galna .
du är uppenbarligen sjuk .
du har slut på ursäkter .
ni har slut på ursäkter .
du har förmodligen rätt .
du är antagligen trött .
ni är antagligen trötta .
du är helt värdelös .
du är för aggressiv .
ni är för aggressiva .
du är väldigt vacker .
din tid är nästan slut .
er tid är nästan slut .
alla vägar leder till Rom .
låt oss sköta vårt jobb .
Tydligen är jag adopterad .
är de här bananerna mogna ?
är du Toms dotter ?
följer någon efter dig ?
kommer ni med oss ?
kommer du med oss ?
är du rädd än ?
är ni rädda än ?
är du bra på tennis ?
är du på biblioteket ?
Hotar ni mig ?
bättre sent än aldrig .
Chefer är också människor .
ring mig när det är färdigt .
ring dem i kväll .
kan jag hämta er någonting ?
kan jag hämta dig någonting ?
kan någon verifiera det ?
kan någon intyga det ?
kan något bekräfta det ?
kan någon bestyrka det ?
kan någon bevisa riktigheten av det ?
kan du vakta ungarna ?
kan du passa barnen ?
kan ni passa barnen ?
kom när du vill .
hände det verkligen ?
hittade dom någonting ?
hittade de någonting ?
tyckte du om matchen ?
hade du roligt på matchen ?
tyckte du om föreställningen ?
hade du roligt på föreställningen ?
tyckte du om rundturen ?
tyckte du om rundvandringen ?
åt du frukost ?
åt ni frukost ?
har du ätit frukost ?
har ni ätit frukost ?
hörde du klickljudet ?
såg du matchen ?
vann du trofén ?
sade jag inte just det ?
drömmer du på franska ?
har du någon lösning ?
har ni någon lösning ?
kan du någon franska ?
vet du vem han var ?
vet ni vem han var ?
tycker du om vitt vin ?
läser du Toms blogg ?
studerar du kemi ?
pluggar du kemi ?
Pluggaru kemi ?
har Tom några söner ?
vet Tom vem jag är ?
ser Tom förvirrad ut ?
blir du ledsen av det ?
gör det dig ledsen ?
gör det er ledsna ?
blir ni ledsna av det ?
var inte fräck emot mig .
Smickra inte dig själv .
lova att du inte blir arg .
få mig inte att skada dig .
få mig inte att döda dig .
få mig inte att döda er .
öppna inte lådan än .
ta inga risker .
berätta inte för din mamma .
slösa inte bort Toms tid .
slösa inte Toms tid .
oroa dig inte . det är enkelt .
oroa dig inte . det är lätt .
Alver har spetsiga öron .
allt är möjligt .
eld är väldigt farligt .
tar du dörren ?
ge mig mikrofonen .
gå hem . vila upp dig .
har du ätit frukost ?
han blåste ut ljuset .
han har inte hatt på sig .
han tycker inte om kaffe .
han är alltid på väg någonstans .
han hoppade över diket .
han levde ett enkelt liv .
han låtsas vara döv .
han kommer nog inte .
han svalde sin stolthet .
han tog fram några mynt .
han tog ut några mynt .
han gör inte en fluga förnär .
han är mörk och snygg .
hennes klänning såg billig ut .
här kommer vår lärare .
historien upprepar sig .
vad sägs om en kopp te ?
hur mycket kostade den där ?
hur mycket är den här värd ?
hur var din dag idag ?
jag råder dig att inte åka .
jag uppskattar din tid .
jag uppskattar ditt jobb .
jag uppskattar ditt arbete .
jag uppskattar ert arbete .
jag tror han är ärlig .
jag tror att han är ärlig .
jag köpte en ny handväska .
jag mutade polisen .
jag kom hit tillsammans med mina vänner .
jag kan inte komma just nu .
jag kan inte hantera det här .
jag kan inte göra det där heller .
jag kan inte gå till polisen .
jag kan inte bara stanna här .
jag kan inte riktigt göra det .
jag kan inte se någonting .
jag kunde inte se någonting alls .
jag köpte inget bröd .
jag köpte inte den där boken .
jag har ingen cykel .
jag gillar inte den här boken .
jag gillar inte ditt namn .
jag vet inte riktigt än .
jag pratar inte japanska .
jag kan inte japanska .
jag förstår mig inte på konst .
jag förstår dig inte .
jag vill inte ha någon frukt .
jag drack igen för mycket .
jag drömde att jag flög .
jag kände mig som ett stort fån .
jag hittade min borttappade plånbok .
jag fick A på min uppsats .
jag antar att Tom inte är hemma .
jag hatar folk som Tom .
jag hatar människor som Tom .
jag hatar personer som Tom .
jag har en katt och en hund .
jag har ett tillkännagivande .
jag har en kungörelse .
jag har ett meddelande .
jag har gjort ett bra jobb .
jag har massor med vänner .
jag måste göra det själv .
jag måste lära mig franska .
jag hör ett konstigt ljud .
jag hörde någon skrika .
jag hörde dörren stängas .
jag hjälpte honom igår .
jag gömde den i min frysbox .
jag hoppas att det inte är sant .
jag hoppas att det där inte är sant .
jag kunde bara inte säga nej .
jag vill bara gå hem .
jag vill bara åka hem .
jag vet knappt någonting alls .
jag vet vad som dödade Tom .
jag bor i en lägenhet .
jag bor i lägenhet .
jag älskar den restaurangen .
jag behöver en extra kudde .
jag behöver lära mig franska .
jag äter bara koscher mat .
jag var bara där en gång .
jag gick bara dit en gång .
jag beställde kinesisk mat .
jag beställde kinesiskt .
jag fick ett jobberbjudande .
jag minns många saker .
jag sa att Tom är en vän .
jag borde vila mig lite .
jag borde få mig lite vila .
jag talar för alla människor .
jag misstänker att Tom är spion .
jag lärde mig franska på egen hand .
jag tycker att Tom är dåraktig .
jag tror att Tom ljög för oss .
jag tycker att han är skicklig .
jag trodde att jag förlorat dig ,
jag trodde att jag förlorat er .
jag trodde att Tom hade stuckit .
jag trodde Tom var död .
jag trodde att du gillade mig .
jag trodde du gillade mig .
jag trodde att ni gillade mig .
jag trodde ni gillade mig .
jag trodde att du tyckte om mig .
jag trodde du tyckte om mig .
jag trodde att ni tyckte om mig .
jag trodde ni tyckte om mig .
jag trodde att du var Tom .
jag tog med mig min kamera .
jag värdesätter vår vänskap .
jag vill göra det själv .
jag vill studera utomlands .
jag vill plugga utomlands .
jag ville rädda dig .
jag var i bergen .
jag var inte det minsta rädd .
jag åkte till sjukhuset .
jag kommer alltid att älska dig .
jag kommer alltid att älska er .
jag hjälper dig gärna .
jag skulle vilja hyra en bil .
jag ringer dig vid sju .
jag hälsar på dig någon gång .
jag är allergisk mot gluten .
jag är glad att vi är överens .
jag går till butiken .
jag har laktosintolerans .
jag bor i stan .
jag letar efter min nyckel .
jag är ingen nybörjare längre .
jag kommer inte att följa med dig .
jag gör bara min plikt .
jag använder datorn .
jag diskar .
jag har alltid haft tur .
jag har bara sett det en gång .
jag har bara sett den en gång .
är någon frånvarande idag ?
är det okej om jag sitter här ?
är det okej om jag sätter mig här ?
går det bra att jag sitter här ?
går det bra att jag sätter mig här ?
finns det vatten på Mars ?
är din mor hemma ?
det är svårt för mig .
den ser ut som en kaktus .
det måste vara skrämmande .
det var extremt roligt .
snart är det vår .
det är en present till dig .
det är en svår situation .
det är nästan omöjligt .
det är alltid mörkt där .
det är närapå omöjligt .
bara följ ditt hjärta .
kom ned från scenen bara .
håll dig undan från hunden .
håll dina händer borta från mig .
skratt smittar av sig .
vi tar det en gång till .
Ligg på din högra sida .
kärleken kommer så småningom .
som tur är blev ingen blöt .
fatta ditt eget beslut .
Mary gillar att titta på tv .
får jag gå på toaletten ?
kan jag få se på matsedeln ?
kan jag få se på menyn ?
Tom kanske kan hjälpa oss .
det mesta är på franska .
mitt skägg växer snabbt .
det värker i hela kroppen .
jag har ont i hela kroppen .
min mamma lagar mat åt mig .
Ljug aldrig igen .
New York är en stor stad .
Pandor är väldigt smarta .
stanna gärna och ät middag .
se saker som de är .
vi ses igen imorgon .
ska jag stänga dörren ?
hon bet i äpplet .
hon är van vid att sitta .
hon vill verkligen gå .
hon har tappat bort bilnyckeln .
hon spelar Monopol .
visa hur man gör det där .
spindlar är inte insekter .
sluta vara så dramatisk .
sluta att bita på naglarna .
sluta bita på naglarna .
säg att du skämtar !
den där kostade mig en förmögenhet .
den där mannen är panikslagen .
kriget tog slut 1954 .
det hade varit roligt .
Publiken applåderade .
Bullen var halväten .
katten satt på mattan .
hunden skrämde katten .
dörren öppnades långsamt .
första gången är gratis .
ju förr desto bättre .
tåget beräknas ankomma kl. 6 .
det var ingen där .
det finns ingen hastighetsbegränsning .
de här är mycket ömtåliga .
de här är väldigt sköra .
de utgör ett skickligt lag .
de säger att kärleken är blind .
de reste tillsammans .
den här konstnären dog ung .
det är ett fritt land .
det här är min väckarklocka .
detta är min vän Tom .
det här är inte en mening .
detta är inte acceptabelt .
den här tidningen är gratis .
den här vägen är farlig .
idag är det den 1 september .
Tom tackade ja till erbjudandet .
Tom har alltid på sig hatt .
Tom bär alltid hatt .
Tom och jag var vänner .
Tom bakade lite muffins .
Tom knäppte sin skjorta .
Tom undanhöll bevis .
Tom kunde tala franska .
Tom kunde inte hitta Mary .
Tom kunde inte finna Mary .
Tom talade inte till mig .
Tom dricker inte så mycket .
Tom dök in i simbassängen .
Tom fritog gisslan .
Tom gav Mary en banan .
Tom har händerna fulla .
Tom har gått ned nästan 14 kilo .
Tom har inget perspektiv .
Tom är granne till Mary .
Tom håller på att bli ursinnig .
Tom håller i en kniv .
Tom är på sjukhuset .
Tom är på väg hit .
Tom är ganska glömsk .
Tom är fortfarande min vän .
Tom är fortfarande skeptisk .
Tom har någonting på gång .
Tom är väldigt rädd .
Tom väntar på dig .
Tom väntar på er .
Tom är inte här längre .
Tom vet att vi litar på honom .
Tom lever ett stillsamt liv .
Tom gjorde många misstag .
Tom begick många misstag .
Tom hade aldrig en chans .
Tom hade aldrig någon chans .
Tom har sällan på sig hatt .
Tom bär sällan hatt .
Tom sa att han är kanadensare .
Tom säger att han inte kommer att rösta .
Tom säger att han är kanadensare .
Tom verkar sova .
Tom har sällan på sig hatt .
Tom bär sällan hatt .
Tom sköt mig i benet .
Tom sov på golvet .
Tom luktade på blomman .
Tom tog av sig skjortan .
Tom tog av sig tröjan .
Tom försökte behålla lugnet .
Tom ville träffa Mary .
Tom föddes på ett skepp .
Tom är för tidigt född .
Tom var min bästa vän .
Tom torkade sig i pannan .
Transplantationer räddar liv .
vi tar kreditkort .
vi har ingen mat .
vi har mycket mat .
vi har inte börjat än .
vi behöver lite mera mat .
vi hyrde en lägenhet .
vi värdesätter våra kunder .
vi vill ha hälsosammare mat .
vi vill ha mer hälsosam mat .
vi planterade träd .
då är det bäst att vi skyndar oss .
vi kommer att överleva .
jag måste bege mig nu .
jag måste ge mig av nu .
vilken fantastisk blomma !
vad är du rädd för ?
vad är ni rädda för ?
vad har vi för val ?
vad tycker du , Tom ?
vad mer behöver repareras ?
vad letade jag efter ?
vad var det du drack ?
vad ska du säga till Tom ?
vad heter Tom i efternamn ?
vad är alternativet ?
vad är det för fel med det ?
vad hette du nu igen ?
vad var det du heter nu igen ?
när kan vi mötas igen ?
när kan vi träffas igen ?
när kan vi ses igen ?
när börjar våren ?
var är Toms saker ?
var är bilnycklarna ?
var kan jag köpa frimärken ?
var kom den ifrån ?
var kom det ifrån ?
var hittade du Tom ?
var fann du Tom ?
var fick du tag på den där ?
vem arbetar vi för ?
vem jobbar vi för ?
vem ska du gå med ?
Vilka ska du gå med ?
vem går du med ?
Vilka går du med ?
vem ska du dit med ?
Vilka ska du dit med ?
vem är du där med ?
vem dansade Tom med ?
vem upptäckte Amerika ?
vem är vi skyldiga pengar ?
Vilka är vi skyldiga pengar ?
vem uppfann pianot ?
vem skulle du rösta på ?
vems resväska är det där ?
vad viskar ni för ?
varför kommer du så tidigt ?
varför ge dem någonting ?
varför var Tom rädd ?
varför frågar du det ?
varför skulle du fråga det ?
kommer Tom att vara här idag ?
i går var det torsdag .
du är längre än mig .
du är längre än jag .
du kan inte gå ut dit .
du får inte gå ut dit .
man kan inte leva för evigt .
du kan inte få oss att sluta .
du kan inte lita på någon .
ni är farliga .
du har ett bra minne .
ni måste ha tålamod .
du ser ut som en apa .
du får inte röka här .
du borde inte vara arg .
du borde inte äta här .
du låter besviken .
ni låter besvikna .
mig lurade du allt .
du skrattar alltid .
du är smartare än jag .
det blåste en kall vind .
en kopp kaffe , tack .
en ponny är en liten häst .
Alle man , överge skeppet !
hela besättningen , överge skeppet !
är det några frågor ?
är du verkligen kanadensare ?
är det mig du menar ?
är du fortfarande arg på mig ?
är ni fortfarande arga på mig ?
fråga henne vad hon har köpt .
var trevligare mot din syster .
var trevligare mot er syster .
svarta katter betyder otur .
ring mig när du kommer tillbaka .
kan någon annan svara ?
kan du räkna på franska ?
kan du föra ett flygplan ?
kan du inte prata engelska ?
rätta mig om jag har fel .
hjälpte Tom dig verkligen ?
sa någon någonting ?
såg du den på riktigt ?
såg du det på riktigt ?
hittade du din handväska ?
hittade du din börs ?
gör som läkaren sagt .
tar ni det här kortet ?
har du några stearinljus ?
har du några vapen ?
tycker du om blåmögelost ?
gillar du att äta fisk ?
gillar du denna trädgård ?
älskar ni er mor ?
behöver du ett kuvert ?
behöver du ett paraply ?
behöver du paraply ?
pratar du med din hund ?
vill du hänga ?
vill ni hänga ?
vill någon ha en öl ?
Ställ inga frågor .
säg aldrig hennes namn .
ge mig inte den där blicken .
låt inte Tom sitta där .
titta inte in i lådan .
vet du inte vem jag är ?
vet ni inte vem jag är ?
känner du inte igen Tom ?
känner ni inte igen Tom ?
det vet vilket barn som helst .
det vet till och med ett barn .
det vet till och med barn .
allt är jättebilligt .
Avgifterna ska snart gå upp .
ta reda på vad Tom vet .
ta reda på vad Tom vill .
ge mig ett exempel till .
Grekland har många öar .
har du varit en stygg pojke ?
har du varit i Boston ?
har ni varit i Boston ?
har du valt ett ämne ?
har du valt ett tema ?
har du hittat någonting ?
har ni hittat någonting ?
har du hört från Tom ?
har ni hört från Tom ?
har du tappat vettet ?
har du inte bestämt dig än ?
han betedde sig som ett barn .
han uppför sig som ett barn .
han valde dem på måfå .
han gick inte upp tidigt .
han steg inte upp tidigt .
han har bytt namn .
han har inte lyckats än .
han är upptagen hela tiden .
han är angelägen att åka dit .
han är flytande på Engelska .
han har inte på sig en hatt .
han har inte på sig hatt .
han har inte hatt på sig .
han har inte en hatt på sig .
han är lång och stilig .
han gick ut i regnet .
han kommer alltid att älska henne .
så här fungerar det .
Hallå , vad gör du ?
hur löste sig allt ?
hur gick det med allt ?
hur hamnade du här ?
hur hamnade ni här ?
hur kom du in hit ?
hur kom ni in hit ?
hur tog du dig in hit ?
hur tog ni er in hit ?
hur kom du in ?
hur tog du dig in ?
hur tänker du hjälpa till ?
hur tror du att jag känner ?
hur tror ni att jag känner ?
hur tror du att jag känner mig ?
hur tror ni att jag känner mig ?
hur långt är det till Boston ?
hur lång är den där bron ?
hur mycket kostar den här kameran ?
hur är ditt liv som gift ?
hur är ert liv som gifta ?
du äcklar mig .
jag är inte på väg någonstans .
jag antar att du har en bil .
jag antar att du har bil .
jag köpte många böcker .
jag köpte en massa böcker .
jag tror inte mina ögon .
jag kan inte knäcka den här koden .
jag kan inte ändra på vem jag är .
jag kan inte göra det själv .
jag klarar det inte själv .
jag kan inte göra det just nu .
jag kan inte göra det längre .
jag kan inte göra det här längre .
jag kan inte låta dig göra det .
jag kan inte låta er göra det .
jag kan inte riktigt minnas .
jag står inte ut med sjukhus .
jag kan inte stå ut med ljudet .
jag kan inte tänka mig något annat .
jag kunde göra det åt dig .
jag kunde inte somna .
jag menade inte något av det .
jag behövde inte din hjälp .
jag behövde inte er hjälp .
jag rörde ingenting .
jag skrev ingenting .
jag skrev inte någonting .
jag känner mig inte särskilt lycklig .
jag måste inte vara här .
jag känner henne inte alls .
jag gillar inte den affären .
jag tycker inte om den affären .
jag tycker inte om det här godiset .
jag tycker om inte den här platsen .
jag gillar inte den här platsen .
jag tycker inte om det här stället .
jag gillar inte det här stället .
jag ser inga blåmärken .
jag vill inte vara rik .
jag vill inte växa upp .
jag vill inte bli vuxen .
jag njuter av klassisk musik .
jag har lust att vara ensam .
jag känner för att vara ensam .
jag tyckte synd om pojken .
jag fick ett F i kemi .
det är nog dags att dra .
jag drömde om honom .
jag har massor av kameror .
jag har en till fråga .
jag har en annan fråga .
jag har en fråga till .
jag har familj i Boston .
jag måste göra det här själv .
jag måste göra detta själv .
jag måste stryka min skjorta .
jag klippte nyss naglarna .
jag tjänade precis tre lax .
jag behöver bara hitta Tom .
jag vill bara ha roligt .
jag vill bara ha kul .
jag vill bara hjälpa er .
jag vill bara hjälpa dig .
jag vet att jag kommer att dö .
jag vet vad det heter .
jag vet vad det kallas .
jag vet att du måste ha fullt upp .
jag vet att du har haft fullt upp .
jag vet att du har varit upptagen .
jag gillar ditt sätt att prata på .
jag gillar hur du pratar .
jag gillar ditt sätt att tala på .
jag gillar hur du talar .
jag tycker om ditt sätt att prata på .
jag tycker om ditt sätt att tala på .
jag tycker om hur du talar .
jag tycker om hur du pratar .
jag tycker om att läsa nyheterna .
jag låste dörren på framsidan .
jag förlorade allt jag hade .
jag förlorade allt som jag hade .
jag gick vilse i Boston .
jag gjorde bröllopstårtan .
jag fattar mina egna beslut .
jag såg det faktiskt aldrig .
jag spelar ofta volleyboll .
jag föredrar cola framför kaffe .
det tror jag verkligen inte .
jag gillar verkligen den där tjejen .
jag gillar verkligen den här boken .
jag behöver verkligen pengarna .
jag behöver verkligen din hjälp .
jag behöver verkligen er hjälp .
jag återvände till huset .
jag cyklade enhjuling idag .
jag sade att det var okej .
jag såg bilen köra på en man .
jag borde inte ha ringt .
jag tror fortfarande på kärleken .
jag känner mig fortfarande inte säker .
jag sträckte ut armarna .
jag sträckte ut benen .
jag behövde plötsligt en bil .
jag antar att du har rätt .
jag tror att jag är utarbetad .
jag tror att jag är överansträngd .
jag tror att jag missade min buss .
jag tycker att Tom är envis .
jag tror att han heter Tom .
jag tror att det är bäst att du går .
jag trodde att jag hörde musik .
jag trodde att jag såg ett spöke .
jag trodde att jag var i tid .
jag trodde att Tom erkände .
jag trodde att alla visste .
jag trodde att vi kunde prata .
jag trodde att du hatade Tom .
jag trodde att du gillade Tom .
jag trodde att du tyckte om Tom .
jag trodde att du åkte hem .
jag trodde att ni åkte hem .
jag trodde att ni gick hem .
jag trodde att du skulle gilla det .
jag trodde att du skulle gilla den .
jag trodde att du skulle tycka om det .
jag trodde att du skulle tycka om den .
jag trodde att ni skulle gilla den .
jag trodde att ni skulle gilla det .
jag trodde att ni skulle tycka om den .
jag trodde att ni skulle tycka om det .
jag sa åt Tom att ta det lugnt .
jag tog en tur till Boston .
jag besökte Tom i Boston .
jag vill ha ett par handskar .
ja vill äta glass .
jag vill äta glass .
jag vill bo i Italien .
jag var inte redo för det här .
jag var inte särskilt nervös .
jag önskar att jag hade vetat .
jag önskar att vi kunde göra det .
jag önskar att vi hade mer tid .
jag undrar om Tom är upptagen .
jag skulle hjälpa dig om jag kunde .
jag skulle hjälpa er om jag kunde .
jag skulle vilja tro dig .
jag skulle vilja tro er .
jag skulle vilja låna den här .
jag skulle vilja låna detta .
jag skulle vilja gå hem nu .
jag skulle vilja betala kontant .
jag skulle vilja träffa Tom nu .
jag skulle vilja sjunga en sång .
jag skulle vilja prata med Tom .
jag skulle vilja tala med Tom .
jag tar det här paraplyet .
jag ska precis äta lunch .
jag är faktiskt väldigt lycklig .
jag kommer till hotellet .
jag är orolig för Tom .
jag ser mig bara omkring .
jag är ganska trött idag .
jag letar efter mina nycklar .
jag gömmer ingenting .
jag döljer ingenting .
jag hemlighåller ingenting .
jag är på åttonde våningen .
jag är stolt över er alla .
jag är stolt över er .
jag har glömt bort hennes namn .
jag har glömt bort hans namn .
jag har hittat en lägenhet .
jag har aldrig hört talas om dig .
du kan gå om du vill .
ni kan gå om ni vill .
är allt under kontroll ?
är det där allt du hade med dig ?
är det här verkligen din bil ?
den verkar vara sönder .
den verkar vara trasig .
det verkar vara brutet .
det gör inte så ont .
det var inte roligt alls .
det är roligt att spela tennis .
det är regn på väg .
det är inte lönt att klaga .
det är rätt beslut .
köp lite godis åt Tom bara .
köp lite godis åt Tom nu .
ta bara ett djupt andetag .
sparka så hårt som du kan .
låt mig ge dig mitt kort .
som jag sa , jag var upptagen .
se på alla dessa lådor .
kan jag använda telefonen ?
Apor är intelligenta .
min bror är lärare .
mitt namn är inte viktigt .
vad jag heter är inte viktigt .
mina föräldrar är skilda .
ingen står över lagen .
ingen av oss talar franska .
det är inte söndag varje dag .
visst , jag förstår .
det är roligt att spela baseball .
Skorpioner är farliga .
hon nickade till svar .
hon gillar inte fotboll .
hon sover redan .
hon kommer kanske i morgon .
hon sa att hon hade en förkylning .
hon hade ont i hela kroppen .
hon gör inte en fluga förnär .
Skriv under på den prickade linjen .
någon förstörde min kamera .
någon gjorde sönder min kamera .
någon hade sönder min kamera .
ta Tom till stationen .
det gäller honom också .
det gäller även honom .
det stör inte Tom .
det där är varför han blev arg .
barnet slutade gråta .
lådan är nästan tom .
lådan var nästan full .
katten fångade råttorna .
katten ligger på bordet .
Kakburken är tom .
hunden är på stolen .
dörren öppnas nu .
Hönan har värpt ett ägg .
Timvisaren är sönder .
huset är sålt .
huset har sålts .
tangentbordet är bakgrundsbelyst .
Damen är över åttio .
flygplanet är överbokat .
Ormen frestade Eva .
Signalen blev grön .
Ormen ömsade skinn .
gatorna är översvämmade .
telefonen är trasig .
de två männen skakade hand .
de två männen tog i hand .
vattnet frös till is .
yoghurten är jättegod .
vad är problemet i så fall ?
det finns inga droger här .
det saknas en gaffel .
det fattas en sida .
det finns en hållplats här .
det finns en busshållplats här .
det finns ett vykort här .
det finns en smörgås här .
det är en smörgås här .
de här skorna passar på mina fötter .
de är korta och smala .
de gick in i djungeln .
de skrattade åt min idé .
de kan gå imorgon .
de erbjöd assistans .
de erbjöd hjälp .
de låter besvikna .
Tänk på din framtid .
den här boken tillhör mig .
den här kon är inte brännmärkt .
den här maten luktar ruttet .
detta är en japansk docka .
det här är en gammal byggnad .
det här kommer att bli roligt .
det var så här det hände .
det här är ganska exakt .
det här är biljettkön .
detta var en skön känsla .
det här var en skön känsla .
Tom gillar faktiskt Mary .
Tom och jag är väldigt upptagna .
Tom bad mig titta förbi .
Tom åt en tidig middag .
Tom tror på älvor .
Tom blåste ut ljuset .
Tom kom tillbaka till Boston .
Tom kan visa dig runt .
Tom kan inte lämnas ensam .
Tom kan inte sjunga höga A .
Tom kan inte sjunga ett högt A .
Tom kan inte arbeta i morgon .
Tom är verkligen snål .
Tom är sannerligen snål .
Tom gjorde det för skojs skull .
Tom dödade ingen .
Tom dödade inte någon .
Tom begick inte självmord .
Tom nämnde inte Mary .
Tom nämnde inte det .
Tom litade inte på någon .
Tom tycker inte om Boston .
Tom behöver ingen käpp .
Tom somnade till slut .
Tom flög hem till Boston .
Tom glömde köpa bröd .
Tom glömde att köpa bröd .
Tom åker till jobbet med bil .
Tom åkte fast för fortkörning .
Tom hade mer arbete att uträtta .
Tom gav asken till Mary .
Tom gav lådan till Mary .
Tom har gjort allt han kan .
Tom har aldrig haft ett jobb .
Tom satte av mot dörren .
Tom är väldigt modig .
Tom är säkert rädd .
Tom är säkert rädd .
Tom håller på att äta frukost .
Tom är trogen Mary .
Tom är Mary trogen .
Tom kommer att klara sig .
Tom döljer någonting .
Tom är maktlysten .
Tom har makthunger .
Tom är makthungrig .
Tom är i nöjesbranschen .
Tom lär sig engelska .
Tom saknar ett finger .
Tom är min storebror .
Tom har timlön .
Tom är mycket fotogenisk .
Tom är blyg och feg .
det var Tom jag ringde .
Tom är väldigt intelligent .
Tom väntar på Mary .
Tom är inte rädd för dig .
Tom är inte bra på att ljuga .
Tom har inte på sig några skor .
Tom stirrade bara på Mary .
Tom vet var Mary är .
Tom tycker om att spela kort .
Tom tittade på sin klocka .
Tom kollade på sin klocka .
Tom tittade på klockan .
Tom kollade på klockan .
Tom tittade på golvet .
Tom tittade i golvet .
Tom tittade in i lådan .
Tom lyssnar aldrig på mig .
Tom öppnade sin resväska .
Tom skalade potatis .
Tom tog upp telefonen .
Tom tycker verkligen om Boston .
Tom sade nästan ingenting .
Tom verkar vara en idiot .
Tom visade Mary lådan .
Tom visade lådan för Mary .
Tom visade asken för Mary .
Tom låter besviken .
Tom tror att han vet varför .
Tom sa att han var upptagen .
Tom brukade köra buss .
Tom var med mig hela dagen .
Tom åkte tillbaka till Boston .
Tom gör inte en fluga förnär .
Tom vred ur trasan .
Tom ! vad sysslar du med ?
Tom ! vad gör du ?
Tom ! vad håller du på med ?
försök att inte äta för mycket .
var någon annan frånvarande ?
vi har alla våra hemligheter .
vi kommer alla att dö .
vi äter frukost .
vi ska mötas vid sju .
vi frågade Tom om det .
vi diskuterade vad vi skulle göra .
vi vill inte avbryta .
vi har tre flygplan .
vi har varit uppe hela natten .
vilken färg har ditt hår ?
vad menar du egentligen ?
vad vill du köpa ?
vad står &quot; PTA &quot; för ?
vad hände i Boston ?
vad är din blodgrupp ?
vad höll Tom på med här ?
vad var det inne i lådan ?
vad gör du idag ?
vad gör du i dag ?
vad väntar du på ?
vad har du för nationalitet ?
när kom han hit ?
när anlände han ?
var är dina bröder ?
var är era barn ?
var kan jag få tag på kartan ?
var var den svarta katten ?
vem håller du på ?
vem hejar du på ?
Vilka håller du på ?
Vilka hejar du på ?
vem väntar du på ?
vem åt den sista kakan ?
varför beskyller du mig ?
varför är du arg på mig ?
varför är du så arrogant ?
varför gick du inte först ?
varför gick ni inte först ?
varför lagar du aldrig mat ?
kan du sätta på teven ?
kan du sätta på tv:n ?
du gjorde ett väldigt bra jobb .
du har inget val .
du ser inte så värst upptagen ut .
du tappade din penna .
du tappade din blyertspenna .
du har ett meddelande här .
du måste låta mig hjälpa till .
du har för mycket att göra .
ni har för mycket att göra .
du är skyldig mig trettio spänn .
du sade att jag skulle bli bättre .
du verkar ganska säker .
ni verkar ganska säkra .
du borde inte tjuvlyssna .
ni borde inte tjuvlyssna .
du tänker på allt .
ni tänker på allt .
du borde inte gå ut .
du är en vacker flicka .
du är en vacker tjej .
ni har helt rätt .
du äger en bil , eller hur ?
du har bil , va ?
ni har bil , va ?
dina gäster väntar .
din önskan har gått i uppfyllelse .
är det någonting jag har missat ?
talar de franska ?
är du lika uttråkad som jag ?
kommer du eller inte ?
är du helt galen ?
är du här tillsammans med någon ?
är du inte klok ?
försöker du fly ?
båda mina fötter är uppsvullna .
bröd är gjort på vete .
hämta lite kallvatten till mig .
hämta mig lite kallvatten .
förresten , var är Tom ?
ring brandkåren !
kan jag avboka den här biljetten ?
kan jag använda din telefon ?
kan du hjälpa mig lite ?
kan du hålla det en hemlighet ?
kom igen , blunda .
nyfiken i en strut .
nyfiken i en strut !
Tandvård är dyrt .
avbröt jag någonting ?
såg du verkligen Tom ?
har du borstat tänderna ?
köpte du medicinen ?
köpte ni medicinen ?
matade du papegojorna ?
sa du att du skulle gå ?
Sydde du den här för hand ?
måste jag göra någonting ?
har vi något annat ?
gör vad han än säger till dig .
kommer du och Tom bra överens ?
får ni många besökare ?
minns ni Tom ?
kommer ni ihåg Tom ?
har du en ordbok ?
har du ett gem ?
har ni några syskon ?
vet du var vi är ?
vet ni var vi är ?
säljer ni väckarklockor ?
hatar du fortfarande franska ?
tror du att jag skämtar ?
tror ni att jag skämtar ?
vet Tom var jag är ?
betyder det att du går med på det ?
betyder det att du håller med ?
be mig inte att inte sjunga
drick inte så mycket öl .
glöm inte att berätta för Tom .
ge inte Tom några idéer .
låt inte Tom spela piano .
låt inte Tom stanna där .
titta inte på kameran .
titta inte in i kameran .
ta det inte personligt .
kasta inte in handduken .
rita en linje med linjal .
kvällen närmade sig .
alla satte sig ner för att äta .
alla pratade om det .
allt var väldigt bra .
fyll burkarna med vatten .
först till kvarn får först mala .
Mjöl är gjort på vete .
ge mig en flaska vin .
morfar köpte den till mig .
ha en underbar kväll .
ha en fantastisk kväll .
har du bestämt dig redan ?
har du någonsin varit på TV ?
har du matat hunden än ?
han erkände sina misstag .
han kom för sent som vanligt .
han kan inte fatta ett beslut .
han har ingen biljett .
han tycker om att spela tennis .
han går i tionde klass .
han tycker mycket om musik .
han låter den här pistolen vara laddad .
han känner många människor .
han lyfte upp henne i luften .
han tycker mycket om musik .
han slutade aldrig att skriva .
han pratade aldrig om det .
han stal plånboken av mig .
han stack sitt hus i brand .
han satte eld på sitt hus .
han lärde sig själv franska .
han kommer vanligtvis i tid .
han brukar komma i tid .
han valdes till president .
han blev ditsatt för mord .
han blev falskeligen anklagad för mord .
han blev snärjd för mord .
han hade snö upp till knäna .
han låg på rygg .
han kommer att älska henne för alltid .
hjälp mig lyfta paketet .
hennes engelska är utmärkt .
hans kropp hittades aldrig .
hans brev gjorde mig arg .
hans tal var för kort .
hur kan ni inte gilla honom ?
hur kan ni inte tycka om honom ?
hur kan du inte gilla honom ?
hur kan du inte tycka om honom ?
hur blir vi av med Tom ?
hur smakar den här soppan ?
hur mycket tycker du om Tom ?
hur mycket gillar du Tom ?
jag är älskad av mina föräldrar .
jag är inte det minsta romantisk .
jag är inte alls romantisk .
jag målar garaget .
jag frågade honom vad han hette .
jag kan inte fatta att jag glömde det .
jag hittar inte det jag vill ha .
jag kan inte gå någon annanstans .
jag minns inte exakt .
jag högg ner ett körsbärsträd .
jag förtjänar en förklaring .
jag gjorde det för tre år sedan .
jag drack inte vattnet .
jag hann inte .
jag ville inte gå hem .
jag tror inte på magi .
jag känner inte för det just nu .
jag mår inte alls bra .
jag känner inte Tom längre .
jag gillar inte modern jazz .
jag tycker inte om det heller .
jag tycker inte alls om det här .
jag gillar inte att titta på tv .
jag tycker inte om dig längre .
jag litar inte på dig heller .
jag har lust att leka med .
jag har också lust att leka .
jag har lust att spela med .
jag har också lust att spela .
jag känner för att spela med .
jag känner för att leka med .
jag känner också för att leka .
jag känner också för att spela .
jag glömde min egen födelsedag .
jag steg upp tidigt i går .
jag växte upp på landet .
jag antar att vi borde gå nu .
jag hade en ordentlig frukost
jag hade ingen aning om vad jag skulle göra .
jag hade ingen aning om hur jag skulle ta mig till .
jag var tvungen att överge min plan .
jag var tvungen att ljuga för alla .
jag var tvungen att fatta ett beslut .
jag har bestämt mig för att gå i pension .
jag har aldrig varit utomlands .
jag måste skriva en essä .
jag har inte tvättat håret .
jag fick höra alltihop .
jag hörde någon skrika .
jag hoppas du har kul .
jag behöver bara lite frisk luft .
jag vet att det inte räcker .
jag vet vad du heter .
jag vet att du fortfarande älskar mig .
jag träffade Tom på flygfältet .
jag behöver en bra ordbok .
jag behöver skölja munnen .
jag har faktiskt aldrig träffat Tom .
jag träffar aldrig Tom längre .
jag tycker verkligen om din musik .
jag tycker verkligen om er musik .
jag sa ju att jag skulle komma på det .
jag såg det för tre timmar sedan .
jag går sällan till biblioteket .
jag tror att jag har allt .
jag tror Tom skulle tycka om det .
jag tror att asken är tom .
jag tror att lådan är tom .
jag trodde att det skulle vara lättare .
jag trodde att du skulle bli arg .
jag talade om allt för mamma .
jag berättade allt för mamma .
jag besökte Paris för länge sedan .
jag väntade i tio minuter .
jag går till arbetet varje dag .
jag promenerar till jobbet varje dag .
jag vill åka dit igen .
jag vill gå dit igen .
jag ville få lite frisk luft .
jag ville överraska henne .
jag blev bortförd av utomjordingar .
jag blev bortförd av rymdvarelser .
jag blev kidnappad av rymdvarelser .
jag blev kidnappad av utomjordingar .
jag var så lycklig på den tiden .
jag önskar att jag vore ung igen .
jag önskar att det vore så enkelt .
jag skulle vilja vara ensam .
jag skulle vilja ha ett glas vin .
jag är där om en stund .
jag tar den gula .
jag tänker inte lyssna på dig .
jag är inte beredd att dö än .
jag målar påskägg .
jag studerar konsthistoria .
jag har redan betalat för den .
jag har alltid velat ha en hund .
är museet öppet idag ?
finns det en app för det ?
är den här buren hajsäker ?
den tillhör min bror .
det stinker verkligen härinne .
det visade sig vara sant .
det var en självmordsbombning .
det var faktiskt mitt fel .
det var inga problem alls .
det var så bullrigt därinne .
det var så stimmigt därinne .
det var så högljutt därinne .
det var inte så dyrt .
det hade varit så enkelt .
det kommer ta några sekunder .
det är skräp . Släng det !
det är jättepinsamt .
det är värt kostnaden .
Koko är en gorillahona .
latin är ett dött språk .
låt mig prata med Tom ensam .
kom så tittar vi i garaget .
se upp för ficktjuvar .
Mary är min före detta flickvän .
får jag låna ditt suddgummi ?
min katt hade ihjäl en ekorre .
min katt dödade denna musen .
min katt dödade den här musen .
min katt dödade denna mus .
min vän studerar koreanska .
min åsikt är irrelevant .
min papegoja dog igår .
min mobil dör snart .
ingen gjorde något annat .
ingen gör någonting .
ingen vill dit .
ingen gör någonting .
nu har jag sett allt .
nu är vi tillsammans igen .
det är klart att jag kommer ihåg dig .
absolut , jag håller helt med .
människorna bodde i byar .
kanske vi möts igen .
hjälp mig med det här är du snäll .
var snäll och sätt på dig skorna .
var snäll och tänd lampan .
var snäll och vänta i fem minuter .
sluta bete dig som ett barn .
russin är torkade vindruvor .
Läs etiketten noggrant .
hon har dåligt rykte .
hon såg upp mot himlen .
hon beställde en kopp te .
sextio nya museer öppnade .
tack för dina kommentarer .
det överraskar mig inte .
det ger mig huvudvärk !
det var bara ett år sedan .
det var för tre veckor sedan .
det var för tre år sedan .
det är struntprat !
det är faktiskt inte sant .
det är verkligen överraskande .
boken kostar fyra dollar .
bussen var nästan tom .
bilen står i garaget .
bilen är i garaget .
skrivbordet är av trä .
maten ser god ut .
Damen förblev tyst .
museet är stängt nu .
den gamla ladan brann ner .
den rosa kudden är ren .
Priserna föll plötsligt .
hyran ska betalas imorgon .
rummet har två fönster .
tåget beräknas ankomma klockan tolv .
det finns för många regler .
det är en katt i lådan .
det finns en telefon här .
det är ingenting här ute .
de är lika starka som vi .
de försökte fly .
de gör så åt alla .
de vet inte vem jag är .
de döpte hunden till Shiro .
de gav hunden namnet Shiro .
de var någon annanstans .
de togs till fånga .
de kommer inte att ha en chans .
de är inte alltid där .
de arbetar på övervåningen .
de är på övervåningen och jobbar .
de är på övervåningen och arbetar .
den här bilen drivs av alkohol .
den här bilen går på alkohol .
detta slott är vackert .
den här maten är glutenfri .
det här gräset behöver klippas .
det här är en vän till mig .
det här är hans bil , tror jag .
detta är hans bil , tror jag .
det här är ganska dyrt .
det här är rätt dyrt .
det här är det värsta av allt .
det här är din sista chans .
det här är ingen tävling .
det här är inte roligt längre .
Tom erkände sitt misstag .
Tom förlorade nästan förståndet .
Tom och de andra håller med .
Tom började må bättre .
Tom kom hit för att hjälpa mig .
Tom kom ut ur grottan .
Tom bestämde sig för att läsa juridik .
Tom gjorde som du föreslog .
Tom fattade det inte heller .
Tom fick det inte heller .
Tom öppnade inte ögonen .
Tom tänkte inte på det .
Tom ser inte nervös ut .
Tom hade många fiender .
Tom har en hel del att förklara .
Tom har mycket att förklara .
Tom har ljugit för mig igen .
Tom har försökt allt .
Tom insisterar på att jag kommer ensam .
Tom har stor fallenhet för idrott .
Tom är plastikkirurg .
Tom är en mycket stark man .
Tom är allergisk mot vete .
Tom grälar med Mary .
Tom bråkar med Mary .
Tom är lika stark som jag .
Tom ligger på rygg .
Tom är en av mina vänner .
Tom är kort för sin ålder .
Tom är väldigt entusiastisk .
Tom är yngre än jag .
Tom söker inte asyl .
Tom vet vad som väntar .
Tom åker om några dagar .
Tom stack för länge sedan .
Tom åkte för tio minuter sedan .
Tom åkte för tre timmar sedan .
Tom älskar chokladtårta .
Tom fick det att se så lätt ut .
Tom måste ha slagit i huvudet .
Tom glömmer aldrig ett ansikte .
Tom lekte med sina katter .
Tom är bra på att spela piano .
Tom skyndade hem från jobbet .
Tom vill verkligen hjälpa till .
Tom sa att han kunde laga den .
Tom säger att Mary är förkyld .
Tom borde uppmuntras .
Tom började bli arg .
Tom berättade för Mary om John .
Tom berättade allt för Mary .
Tom stängde av alarmet .
Tom stängde av radion .
Tom knäppte upp sin skjorta .
Tom brukade stiga upp tidigt .
Tom gick in i cellen .
Tom vill ha någonting annat .
Tom vill någonting annat .
Tom kunde inte svara .
Tom ger inte upp så lätt .
Tom undrar om det är sant .
Skruva ned tv:n .
vi är benägna att slösa tid .
vi gör ingenting .
vi kan ta hissen .
vi beställde ingenting .
vi har inte beställt någonting .
vi sysslar inte med det längre .
vi håller inte på med det längre .
vi har mer än tillräckligt .
vi har bara två dollar .
vi har trettio anställda .
vi har inte gjort någonting .
vi måste gå med en gång .
vi var ett perfekt par .
vi klagar alltid .
det gick ju smärtfritt .
vad firar ni ?
vad firar du ?
vad antyder du för något ?
vad är det du insinuerar ?
vad är det du antyder ?
vad är det ni antyder ?
vad är det ni insinuerar ?
vad antyder ni för något ?
vad skrattar du åt ?
vad tänker du på ?
vad väntar du på ?
vad ville Tom äta ?
vad menar du med det ?
vad behöver du veta ?
vad behöver ni veta ?
vad betyder det här ordet ?
vad är det här för slags hund ?
vad handlar mötet om ?
när kan jag träffa Tom igen ?
när kan jag se dig igen ?
när gifte du dig ?
vart är du på väg ?
var får jag tag på böcker ?
Vilka är alla de här människorna ?
vem tror du att du är ?
varför följer du efter mig ?
varför förföljer du mig ?
varför förföljer ni mig ?
varför följer ni efter mig ?
varför är du på det här skeppet ?
varför är ni på det här skeppet ?
varför är ni på detta skepp ?
varför är du på detta skepp ?
varför kan vi inte göra om det ?
varför kan vi inte göra det igen ?
varför köpte du en blomma ?
varför köpte du en sköldpadda ?
varför köpte ni en sköldpadda ?
varför köpte du den här bilen ?
varför ser du bekant ut ?
varför är fisk så dyrt ?
varför skulle jag säga någonting ?
varför skulle det vara lättare ?
hinner du ?
utan dig är jag ingenting .
kvinnor tjänar mindre än män .
vill ingen sitta med mig ?
i går var en bra dag .
du fattar inte , eller hur ?
ni fattar inte , eller hur ?
du känner inte mig över huvud taget .
ni känner inte mig över huvud taget .
du fick betalt , eller hur ?
du har ingen aning , eller hur ?
du måste lämna Boston .
du kände Tom , eller hur ?
ni vet att jag älskar er båda .
du vet att jag älskar er båda .
du bor här , eller hur ?
du måste vara Toms far .
du äger en bil , eller hur ?
ni äger en bil , inte sant ?
du sa att det var för lätt .
du sade att det var för lätt .
du sade att det var för enkelt .
du hade rätt hela tiden .
du är smartare än jag .
du är smartare än vad jag är .
du är den bästa pappan någonsin .
din franska är utmärkt .
din dotter går på droger .
all kunskap är inte till godo .
är du höjdrädd ?
kommer du att använda den här ?
är du verkligen så naiv ?
det var i alla fall inte tråkigt .
den delen är i alla fall sann .
den delen är åtminstone sann .
att vara ärlig är svårt .
båda är lärare .
bröd bakas i ugn .
bröd bakas i en ugn .
kan jag köpa enbart linserna ?
får jag använda din ordbok ?
barn tycker om sagor .
kom och drick te med mig .
kunde det vara ett mord ?
skulle du kunna vara tyst , tack ?
sa verkligen Tom det ?
lade du märke till några fel ?
upptäckte du några fel ?
beställde du inte rödvin ?
dinosaurier är nu utdöda .
tror du på älvor ?
har ni Guinness här ?
har du ett kreditkort ?
har ni några frågor ?
tycker du om japansk mat ?
tycker ni om att spela spel ?
behöver ni dricka vin ?
har rummet ett badkar ?
bli inte alltför bekväm .
titta inte ut genom fönstret .
vill du inte se Tom ?
rita ett streck på ditt papper .
alla vet vem Tom är .
Tyskland gränsar till Frankrike .
Häng upp din kappa , tack .
Häng din hatt på kroken .
har du någonsin blivit bestulen ?
har jag inte lidit tillräckligt ?
har jag inte lidit nog ?
har jag inte lidit så det räcker ?
hon åt en bit av tårtan .
han blev en berömd sångare .
han köpte ett par skor .
han högg ner ett körsbärsträd .
han bestämde sig för den röda bilen .
han höll henne i ärmen .
han längtar efter att åka utomlands .
han dagdrömmer jämt .
han är arton månader gammal .
han är antingen full eller tokig .
han bor hos sina föräldrar .
han tillverkade en liten hundkoja .
han måste komma söderifrån .
han stod bakom stolen .
han var mina första pojkvän .
han slipade en kniv .
han tittar på dinosaurier .
hjälp mig en minut bara .
hennes hobby är bodybuilding .
här är mitt körkort .
hans tillstånd är kritiskt .
hur gick din intervju ?
hur gick det på din intervju ?
hur gillar du staden ?
hur många bor här ?
vad kostar en öl ?
hur ofta äter du fisk ?
hur allvarlig är krisen ?
jag är ingen morgonmänniska .
jag frågade Tom vad han menade .
jag tror att han heter Tom .
jag är med i en tennisklubb .
jag hittar inte den inställningen .
jag kan inte gå förrän han kommer .
jag kan inte låta dem fånga mig .
jag minns ingenting .
jag kommer inte ihåg vad hon heter .
jag minns inte hennes namn .
jag vill inte ha era hus .
jag vill inte ha dina hus .
jag har inga bröder .
jag har inte tid att laga mat .
jag har inte tid att läsa .
jag förstår det inte heller .
jag vill inte ha någon annan .
jag tvivlar på att Tom är glad .
jag tvivlar på att Tom är lycklig .
jag fick reda på var hon var .
jag har en vän vid namn Tom .
jag har en överraskning åt dig .
jag har en överraskning åt er .
jag har en ätstörning .
jag har lånat två böcker .
jag älskar reor .
jag vet absolut ingenting .
jag behöver myggmedel .
en gång fann jag en bok där .
jag väger bara 45 kilo .
jag spelade fotboll igår .
jag spelade fotboll i går .
jag låtsades arbeta .
jag såg det med mina egna ögon .
jag kommer fortfarande ihåg hans namn .
jag tror att du har rätt .
jag trodde att Tom skulle få panik .
jag trodde att Tom skulle gripas av panik .
jag trodde att Tom skulle råka i panik .
jag trodde att Tom skulle bli panikslagen .
för länge sedan besökte jag Kanada .
jag vill ha tillbaka mina tjugo dollar .
jag vill bli doktor .
jag vill bli läkare .
jag vill att du kommer tillbaka till Boston .
jag var hos en kompis .
jag tittade på tv i morse .
jag önskar att jag hade fler vänner .
jag önskar att alla gillade mig .
jag önskar att alla tyckte om mig .
det skulle jag inte ha gjort .
jag kommer förklara incidenten .
jag är faktiskt ganska trött .
jag är på polisstationen .
jag går ut en stund .
jag går ut ett slag .
jag håller på att lära mig att köra bil .
jag mår inte så bra .
jag ska inte göra illa dig .
jag är inte intresserad av Tom .
jag är ledsen att jag tog upp det .
Förlåt för igår .
Förlåt för i går .
tyvärr , jag har ingen aning .
jag är övertygad om att du är väldigt upptagen .
du är säkert väldigt upptagen .
jag försöker skydda Tom .
jag ser väldigt mycket fram emot det .
jag har aldrig träffat Toms fru .
jag har bara varit där en gång .
jag har sett dig spela tennis .
jag har stängt alla sex fönster .
om du vill prata , prata .
om du vill prata så prata .
om du vill prata , prata då .
Illusioner är kortlivade .
om två dagar fyller jag 13 .
finns det en telefon här ?
är det inte alltid så ?
det blir nog inte lätt .
är inte det vad de vill ha ?
det tar inte särskilt lång tid .
det är lätt att spela tennis .
klockan är sju i London nu .
hon är sju i London nu .
det är deras rätt att rösta .
det är vad alla säger .
det blir troligtvis inte lätt .
det regnade kraftigt hela dagen .
det var bara en tursam gissning .
det var bara början .
det ska bli skönt att komma hem .
det är en svår fråga .
det är mycket mer än så .
det är mycket att tänka på .
den är alldeles underbar .
det är lättare än det ser ut .
det är roligt att spela baseball .
det är skönt att vara hemma igen .
det är mycket enklare såhär .
det är inte en kuggfråga .
det är bara för några veckor .
det gäller bara några veckor .
det är faktiskt inte så mycket .
det är faktiskt väldigt irriterande .
det är dags att gå till skolan .
säg till vad jag kan göra .
låt mig bjuda dig på middag .
låt mig fundera en minut .
Mary gillar mjölk väldigt mycket .
Mary svär som en sjöman .
kan jag få din uppmärksamhet ?
kan jag få er uppmärksamhet ?
min lägenhet är i närheten .
min lägenhet ligger här i närheten .
min hund skäller hela tiden .
min far älskar min mor .
min far är duktig på att simma .
min mamma jobbar på fabrik .
mitt namn står inte med på listan .
min åsikt var irrelevant .
min katt dog i går .
mina planer misslyckades rejält .
mina planer misslyckades kapitalt .
naturen är full av mysterium .
ingen kommer någonsin att få reda på det .
det händer aldrig någonting här .
det är inget fel med Tom .
vänta lite nu .
en kopp kaffe , tack .
vår lärare skrattar sällan .
var snäll och låt Tom göra sitt jobb .
Kavla upp din högerärm .
säkerhet kommer alltid först .
ska jag hålla dig informerad ?
hon skrek till av förvåning .
hon gav mig flera böcker .
hennes arm är gipsad .
hon är ute efter ett bättre jobb .
hon är ingen vanlig sångerska .
borde jag be Tom om ursäkt ?
borde du inte använda handskar ?
någon är i vårt garage .
någon ringde på dörrklockan .
någon stal mitt pass .
fortkörning förorsakar olyckor .
sluta vara så tjurskallig !
tack för rättelsen .
tack för ditt hårda arbete .
tack för ert hårda arbete .
tack så mycket för middagen .
det hände egentligen inte .
det var en lögn , eller hur ?
det skulle inte förvåna mig .
det kommer försätta dig i fara .
det är alldeles korrekt .
det är allt jag behöver för tillfället .
det är käringprat .
Publiken såg uttråkad ut .
lådan var full av böcker .
företaget gick i konkurs .
matchen slutade oavgjort .
matchen blev oavgjord .
mördaren avrättades .
de gamla reglerna gäller inte .
festen spårade ur .
telefonen är trasig .
Posten är stängd .
det är mulet idag .
Soldaten uppgav sitt namn .
tåget har inte kommit ännu .
det finns åtskilliga orsaker .
det har kommit ett brev till dig .
det fanns inte tillräckligt med bränsle .
det finns mycket mer att se .
det finns en restaurang här .
det finns mat på bordet .
det finns ingen plats här .
de här skorna passar perfekt .
de kommer inte idag .
de kan inte heller höra mig .
de byggde en bro .
de steg in i hissen .
de planerar att ordna en fest .
de frös ihjäl .
den här tv:n gjordes i Kina .
den här filmen är sevärd .
det här är en läsvärd bok .
det här är Japans flagga .
den här whiskyn är för stark .
Tom trodde faktiskt på dig .
Tom och jag var båda glada .
Tom kan inte förneka det längre .
Tom samlade på kaffekoppar .
Tom tyckte inte om den idén .
Tom verkar inte hålla med .
Tom gav mig några dollar .
Tom fick en fortkörningsbot .
Tom börjar bli ett problem .
Tom håller på att bli ett problem .
Tom är oerhört upptagen just nu .
Tom är oerhört romantisk .
Tom är muskulös , eller hur ?
Tom är positiv , eller hur ?
Tom är den perfekta pappan .
Tom skickade precis ett mejl till mig .
Tom mejlade mig precis .
Tom skickade precis ett e @-@ postmeddelande till mig .
Tom visste att jag hade rätt .
Tom tycker om att skriva poesi .
Tom gillar att skriva poesi .
Tom behöver kanske inte vår hjälp .
Tom sa att han inte kunde gå .
Tom satt på en närliggande bänk .
Tom säger att det var din idé .
Tom verkar vara väldigt upptagen .
Tom borde ha blivit varnad .
Tom visade Mary pappret .
Tom visade Mary fotot .
Tom smällde igen dörren stängd .
Tom skar av Marys hals .
Tom har ibland på sig en hatt .
Tom har fortfarande mitt paraply .
Tom har mitt paraply fortfarande .
Tom har fortfarande inte dykt up .
Tom ser fortfarande deprimerad ut .
Tom ser fortfarande förvånad ut .
Tom verkar fortfarande bekymrad .
Tom kämpade för att bli fri .
Tom trodde att Mary var upptagen .
Tom sade till Mary att han var upptagen .
Tom sade till mig att den blev stulen .
Tom berättade några snuskiga skämt .
Tom tog av sin gasmask .
Tom försökte väcka Mary .
Tom stängde av apparaten .
Tom fick antibiotika .
Tom var gift på den tiden .
Tom var faktiskt inte där .
Tom har på sig hatt varje dag .
Toms pappa var präst .
Toms mamma dog 2013 .
tänder du lyset ?
vi visste inte vad vi skulle göra .
vi träffas här en gång i månaden .
vi är ingifta släktingar .
vi har alltid varit vänner .
vi har slut på bensin .
vi har slut på fotogen .
vilket stort hus du har !
vilket stort hus ni har !
vad gjorde han efter det ?
vad vill du att jag ska göra ?
vad vill du titta på ?
vad ligger växelkursen på ?
vilken tid passar dig ?
vilken tid passar er ?
vad är klockan i Boston ?
vad var din plan egentligen ?
hur är det att vara döv ?
vad är det för filtillägg ?
vad är filtillägget ?
vad heter den här gatan ?
vad är din fars namn ?
när slutar din lektion ?
när börjar din resa ?
var är de andra flickorna ?
var ligger damernas ?
vart vill du helst åka ?
var ska Tom bo ?
var finns närmaste hotell ?
var ligger närmaste hotell ?
vilket märke gillar du ?
vem målade den här tavlan ?
vem målade den här målningen ?
vem vill ha en bit tårta ?
vem pratade ni med ?
vem pratade du med ?
Vilka pratade du med ?
vad tittar du på mig för ?
vad tittar ni på mig för ?
varför låste du dörren ?
varför trodde du inte på mig ?
varför skrattar alla ?
varför borde jag studera franska ?
varför var Tom inte här idag ?
kommer du göra det med Tom ?
kan du vara snäll och sätta dig ner ?
vill du göra mig sällskap ?
yoga hjälper henne att vara lugn .
du kan inte göra det längre .
du kunde inte kontaktas .
ni kunde inte bli kontaktade .
du behöver inte göra det .
ni behöver inte göra det .
du dricker för mycket kaffe .
du har fel nummer .
du måste göra dina läxor .
du måste återbetala dina skulder .
ni måste återbetala era skulder .
du borde äta mer frukt .
det är bäst att du inte berättar för honom .
det är bäst att ni inte berättar för honom .
en dag kommer du att förstå .
du har alldeles rätt .
du har stavat mitt namn fel .
ni har stavat mitt namn fel .
du har felstavat mitt namn .
ni har felstavat mitt namn .
du har stavat fel på mitt namn .
ni har stavat fel på mitt namn .
en student vill träffa dig .
det är en student som vill träffa dig .
flygplan landar på flygplatser .
allt du behöver göra är att tala .
är jag så olik dig ?
vem som helst kan göra misstag .
arabiska är mitt modersmål .
är mina kläder redan torra ?
ber du om min hjälp ?
kommer du att stanna länge ?
är du redo att beställa nu ?
är ni redo att beställa nu ?
stannar du och äter middag ?
Bankerna öppnar klockan nio .
kan du få ut mig härifrån ?
kan ni få ut mig härifrån ?
kommer du ihåg det här spelet ?
kommer du ihåg den här leken ?
kommer ni ihåg den här leken ?
kommer ni ihåg det här spelet ?
minns du det här spelet ?
minns ni det här spelet ?
kan jag inte stanna här med dig ?
kan du vara lite mer specifik ?
lovade Tom att göra det ?
har allt det här faktiskt hänt ?
läste du verkligen det ?
har du hört vad som hänt ?
har du hört vad som har hänt ?
ser du någonting annat ?
har din mor gjort de där ?
har din mamma gjort de där ?
titta inte ut genom fönstret .
vet de vad som hände ?
säljer de Guinness här ?
vet du vem som dödade Tom ?
tycker du om Ikeamöbler ?
tycker du om de här örhängena ?
gör det något om jag stannar här ?
behöver du någonting annat ?
vill du verkligen hjälpa till ?
vill ni verkligen hjälpa till ?
ångrar du det som du gjorde ?
tror du att Tom var full ?
är det möjligt , tror du ?
är det möjligt , tror ni ?
gör Tom så här varje dag ?
vet Tom att Mary är här ?
öppna inte presenten än .
sätt dig inte på soffan .
sätt er inte på soffan .
rita en bild av dig själv .
alla var väldigt glada .
alla var jätteglada .
Snabbmat kan vara beroendeframkallande .
fyll flaskan med vatten .
ge Tom något att dricka .
Grekerna äter ofta fisk också .
är tåget försenat ?
har du någonsin sett Tom äta ?
har du någonsin sett en val ?
har ni någonsin besökt Rom ?
har du träffat alla här ?
har ni träffat alla här ?
han drog det kortaste strået .
han steg upp klockan fem som vanligt .
han steg upp klockan fem som han brukar .
han har alltid något fuffens för sig .
han är galen i baseboll .
han sitter på stolen .
han lät mig sova över en natt .
han tycker om att vara busig .
han hittade på hela historien .
han såg en hund i närheten av dörren .
han rakade av sig mustaschen .
han talar lite engelska .
han blev attackerad av en haj .
han attackerades av en haj .
han tittade på en svensk film .
han jobbade hårdare än någonsin .
han är lärare , och det är jag med .
han kommer alltid för sent till timmen .
han kommer alltid för sent till lektionen .
han är alltid sen till lektionen .
han tittar alltid på dig .
han läser alltid serietidningar .
han gräver sin egen grav .
han är någonstans i parken .
han är lagkapten .
Nederländerna är ett litet land .
hur fick du in den hit ?
hur fick du in det hit ?
hur har du skadat din hand ?
hur har du tillbringat dagen ?
hur länge sedan hände det ?
hur länge har Tom varit här ?
hur länge har vi varit här ?
hur mycket tid kommer vi att ha på oss .
hur ofta händer det ?
skynda på och ät upp .
jag har alltid velat göra det .
jag antog att det var gratis .
jag antog att den var gratis .
jag har köpt lite aspirin till dig
jag kan inte låta dem fånga dig .
jag kan inte se skillnaden .
jag kan inte stoppa blödningen .
jag skulle behöva lite hjälp här .
jag trodde inte mina ögon .
jag kunde inte låta det hända .
jag kunde inte låta det ske .
jag kunde inte lägga band på mig själv .
jag kunde inte tygla mig själv .
jag kunde inte tygla mig .
jag kunde inte lägga band på mig .
jag ställde inga frågor .
jag bad inte om din hjälp .
jag bad inte om er hjälp .
jag åt ingenting annat .
jag såg ingen som åt .
jag såg inte att någon åt .
jag klandrar dig inte för det här .
jag är inte så förtjust i grönt te .
jag bryr mig inte om vad som hände .
jag går inte ut och äter så ofta .
jag vill inte ens ha dig här .
jag vill inte ens ha er här .
jag har inget val här .
jag har inga lektioner idag .
jag har inga lektioner i dag .
jag känner inga blinda män .
jag vet inte om jag kan hjälpa .
jag gillar inte din attityd .
jag behöver inte mera hjälp .
jag kommer inte ihåg ditt namn .
jag delar inte din åsikt .
jag tror inte att han kommer .
jag vill inte ha mer att dricka .
jag vill inte störa Tom .
jag vill inte bo ensam .
jag tycker om att se på när Tom dansar .
jag känner mig helt hjälplös .
jag känner mig energisk och lycklig .
jag känner mig som en annan person .
jag antog att jag skulle vara säker här .
jag glömde stänga dörren .
jag köpte något att äta till dig .
jag växte upp med att titta på Pokémon .
jag är väl lite full .
det kan väl inte hjälpas .
jag antar att det inte kan hjälpas .
jag har en vän i England .
jag har matteläxa idag .
jag har ingen aning om vem du är .
jag har något i ögat .
jag måste gå på toaletten .
jag hoppas att ni trivs här .
jag hoppas att du trivs här .
jag hoppas att du tycker om att vara här .
jag hoppas att ni tycker om att vara här .
jag tror bara att Tom var full .
jag visste att det inte skulle vara lätt .
jag visste att du kunde svaret .
jag visste att du skulle trivas här .
jag visste att ni skulle trivas här .
jag vet var Tom gömmer sig .
jag gick från festen för tidigt .
jag släppte in katten i mitt rum .
jag tycker mer om katter än hundar .
jag gillar att ha mycket att göra .
jag fick dig att skratta , eller hur ?
jag fick er att skratta , eller hur ?
jag behöver en bättre ordbok .
jag behöver parkera min bil här .
jag måste förnya mitt ID @-@ kort .
jag måste låsa upp den här dörren .
jag behöver din hjälp här .
jag har aldrig menat dig något illa .
jag betalade honom fem dollar .
jag hoppas verkligen att du har rätt .
jag hoppas verkligen att ni har rätt .
jag rev upp kuvertet .
jag sa att jag var förvirrad .
jag sa att det inte var någon här .
jag borde ha studerat flitigare .
jag borde egentligen inte vara här .
jag visade för dem hur man gör .
jag studerar kinesiska i Beijing .
jag tackade Tom för hans hjälp .
jag tror att jag skall köpa en ny bil .
jag tror att jag ska raka huvudet .
jag tror att Tom ville ha min hjälp .
jag tror inte att Tom skulle hålla med .
jag tror hon är 40 år .
jag tror att hon kommer .
jag tror att hon kommer att komma .
jag trodde att jag förstod dig .
jag trodde att det skulle vara värt det .
jag tänkte att det skulle vara värt det .
jag trodde att du var i tjänst .
jag sa till Tom att möta mig här .
jag brukade tycka om att komma hit .
jag bär vanligtvis inte hatt .
jag vill bli taxichaufför .
jag vill förändra världen .
jag vill bo i staden .
jag varnade honom för faran .
jag letade efter min dagbok .
jag satt uppe hela natten och läste .
jag önskar att Tom fortfarande var här .
jag undrar hur det gick till .
kan jag få ett kvitto , tack ?
jag skulle vilja byta rum .
jag skulle vilja byta plats .
jag skulle vilja se dem igen .
jag skulle vilja träffa dem igen .
jag kollar i källaren .
jag är rädd för vilda djur .
jag är medveten om dina problem .
jag är glad att du kunde komma .
jag kommer att sakna er .
jag kommer att sakna dig , Tom .
jag ska ha fest .
jag ska ordna en fest .
jag är glad att du är här , Tom .
jag är i Hong Kong just nu .
jag utreder ett mord .
jag åker om tio minuter .
jag åker på morgonen .
jag ska träffa Tom om en timme .
jag är nära tågstationen .
jag är inte rädd för dig , Tom .
jag är inte tillräckligt erfaren .
jag kommer inte från en rik familj .
jag målar ett påskägg .
jag börjar känna mig trött .
jag säger åt dig att hålla käft .
jag har alltid hatat mörkret .
jag har varit hos tandläkaren .
jag har haft en jobbig eftermiddag .
jag har känt Tom länge .
jag har gjort så många misstag .
jag har börjat röka igen .
faktum var att han till och med älskade henne .
med andra ord : han är lat .
är Tom stor nog att dricka alkohol ?
räcker tiotusen yen ?
är det en seriös fråga ?
är det det som hände här ?
är det vad som hände här ?
ligger hotellet långt härifrån ?
är det långt till hotellet härifrån ?
finns det en busshållplats här i närheten ?
finns det ett apotek i närheten ?
händer detta verkligen ?
äter inte Tom frukost ?
ska inte Tom äta frukost ?
är inte Tom och äter frukost ?
håller inte Tom på och äter frukost ?
håller inte Tom på att äta frukost ?
är inte den där kjolen för kort ?
det snöar nästan aldrig här .
det kan inte ha varit lätt .
jag blev inte klok på det .
jag förstod mig inte på det .
det har snöat i två dagar .
det har inte alltid varit lätt .
det är roligt att spela baseball .
det gjorde mig ytterst glad .
det påverkade egentligen inte oss .
det var faktiskt inte så svårt .
det borde inte ha hänt .
det var ett totalt misslyckande .
det var nästan som en dröm .
det är precis som jag förväntade mig .
det kommer att ta ett tag .
det är inte värt besväret .
det är uppenbart att Tom ljög .
det är antagligen bara ett rykte .
det är faktiskt ganska vanligt .
det är dags för dig att gå .
det är dags att gå till gymmet .
berätta bara vad som hände .
låt oss spela detta spel igen .
långa kjolar är på modet .
Marconi uppfann radion .
Mary är modedesigner .
får jag raka av dina polisonger ?
mjölk är en populär dryck .
min franska håller på att bli rostig .
min franska börjar bli rostig .
jag fyller år i november .
min födelsedag är i november .
min födelsedag är den 22 mars .
min bil står dig till buds .
min framtid ligger i dina händer .
min framtid ligger i era händer .
min farbror är en usel bilförare .
min farbror är usel på att köra bil .
nästa gång ska jag anstränga mig mera .
nästa år blir spännande .
ingen är för gammal för att lära sig .
ingenting kommer att hända .
ingenting sådant hände .
nu ska vi se vad som händer .
Fortsätt med arbetet nu .
ett år består av tolv månader .
Ställ den var som helst .
var snäll och säg åt Tom att vi är här .
vi ses i skolan imorgon .
hon övergav sina barn .
hon kom inte förrän två .
hon kom inte innan två .
hon verkade inte intresserad .
hon talar lite arabiska .
hon nekade mitt önskemål .
hon är gift med en tandläkare .
hon sitter på bänken .
hon börjar irritera mig .
borde jag vänta på Tom här ?
borde vi inte hämta våra saker ?
borde vi inte låsa ?
borde vi inte säga någonting ?
borde du inte ta en paus ?
Rökning är förbjudet här .
det är någon som väntar på dig .
förr eller senare kommer du att ångra det här .
en dag kommer du att ångra det här .
förr eller senare kommer ni att ångra det här .
det är någon som försöker ta sig in .
det är någonting på gång här .
det är någonting lurt på gång här .
det är något som inte stämmer här .
något är inte rätt här .
ta en tupplur om du är trött .
Meddela Tom när du är klar .
berätta för mig hur du känner dig .
säg till när Tom är här .
tack för informationen .
det kommer inte att hända .
det kommer inte att ske .
det var inte det som hände .
det där var en utmärkt putt .
det ska aldrig hända igen .
det är allt jag vet säkert .
det var allt jag ville säga .
det är allt jag har att säga .
det är bättre än ingenting .
det är precis vad jag behöver .
det var precis det jag sa .
det duger åt Tom .
det var precis vad jag behövde .
det är mycket viktigare .
det behövs inte längre .
det angår inte mig .
det är inte svårt att göra .
det kommer inte att bli roligt .
det kommer inte att ske .
så kommer det inte att bli .
det var inte så det gick till .
det är inte mitt problem , Tom .
det är inte därför du är här .
det angår inte mig .
det är en av mina favoriter .
det är bara halva sanningen .
det kommer inte på fråga .
det är precis det det handlar om .
det är antagligen ett tryckfel .
det är orsaken till varför jag är här .
det var så det gick till .
det är otroligt dumt .
det brukar vara ett bra tecken .
det trodde jag också .
det är vad jag har fått höra .
det är vad jag har hört .
det var där Tom och jag träffades .
det var därför vi skilde oss .
tv:n var på hela tiden .
teven var på hela tiden .
Titanic krockade i ett isberg .
väckarklockan ringer .
Skytten dödade hjorten .
Bågskytten dödade hjorten .
boken föll på golvet .
katten klängde vid hennes klänning .
katten är under bordet .
katten ligger under bordet .
staden föll i fiendernas händer .
jag får inte upp skåpdörren .
hunden grävde en grop .
hatten passar henne perfekt .
huset är målat i vitt .
barnen var inte imponerade .
mötet varade till 5 .
den andra fungerar inte .
rummet är fullt av folk .
Ormen svalde en groda .
Teservisen är inte komplett .
tåget är försenat .
det är en stor storm på väg .
taket läcker .
det är absolut riskfritt .
det skadar inte att titta .
det finns ingen orsak till oro .
det finns ingen väg ut härifrån .
det är ingen vid dörren .
det finns ingenting Tom kan göra .
det finns ingenting mer att göra .
det finns ingenting att förklara .
det finns ett litet problem .
det är snö på marken .
det finns så mycket kvar att göra .
det är någon där ute .
det är någonting där inne .
de här ljusen är inte vita .
de här stearinljusen är inte vita .
de behöver inte mig längre .
de behöver mig inte längre .
de serverar inte det här .
det serveras inte här .
de lät mig välja en present .
de betedde sig underligt .
de kommer att heja på er .
de kommer nog på någonting .
de är syskon .
den här boken behandlar Kina .
detta uttryck är arkaiskt .
den här filmen är ett mästerverk .
det här kommer aldrig att ta slut .
det här är inte längre relevant .
det här gör det inte precis bättre .
i morse klarnade det .
det här liknar trakasseri .
det här borde inte vara så svårt .
det här jobbet var svårt att få .
det här ordet kommer från grekiskan .
den här yoghurten smakar konstigt .
de där tulpanerna är vackra .
Tom råkade skjuta Mary .
Tom beundrade Marys mod .
Tom dog nästan den natten .
Tom och Mary blev veganer .
Tom bad Mary att hjälpa honom .
Tom frågade mig vad som hände .
Tom bad oss att följa honom .
Tom bad oss att följa med honom .
Tom köpte en lädersoffa .
Tom köpte en ros åt Mary .
Tom var nära att drunkna .
Tom kom tre timmar för tidigt .
Tom kan köra gaffeltruck .
Tom tycker helt klart om att köra bil .
Tom stängde kontorsdörren .
Tom kunde ha räddat sig själv .
Tom skulle kunna ha rättat sig själv .
Tom skulle kunna räddat sig själv .
Tom gjorde det utan min hjälp .
Tom hittade inte det jag gömde .
Tom hittade inte det som jag gömde .
Tom hittade inte vad jag gömde .
Tom gav mig inga detaljer .
Tom gick inte in på några detaljer .
Tom sa inte vad han gjorde .
Tom verkade inte så glad .
Tom verkade inte så värst glad .
Tom vann inte tävlingen .
Tom dricker inte rödvin .
Tom vet inte vad jag gör .
Tom körde tillbaka till bondgården .
Tom körde tillbaka till farmen .
Tom körde tillbaka till gården .
Tom blinkade med helljusen .
Tom har ofta på sig en hatt .
Tom gav mig trettio dollar .
Tom kom dit före mig .
Tom tog sin examen vid Harvard .
Tom utexaminerades från Harvard .
Tom avlade sin examen vid Harvard .
Tom var tvungen att fatta ett beslut .
Tom har kommit fram till ett beslut .
Tom har druckit en hel del .
Tom har bett om vår hjälp .
Tom började gå mot dörren .
Tom bjöd in Mary till Boston .
Tom är usel på att köra bil .
Tom är skolbusschaufför .
Tom kan köra bil .
Tom är redan ganska full .
Tom är en mycket bra chaufför .
Tom är jättebra på att köra bil .
Tom är i behov av vår hjälp .
Tom gör bara sin plikt .
Tom ligger på backen .
Tom är gammal nog att dricka alkohol .
Tom är ute och går med hunden .
Tom studerar vid Harvard .
Tom borde vara här .
Tom är ofattbart dum .
Tom är väldigt rik , eller hur ?
Tom är väldigt lång , eller hur ?
Tom har på sig en svart hatt .
Tom bär en svart hatt .
Tom sitter och jobbar vid sitt skrivbord .
Tom sitter vid sitt skrivbord och skriver .
Tom är inte Marys pojkvän .
Tom är inte särskilt upptagen , eller hur ?
Tom är väl inte särskilt upptagen ?
Tom är inte särskilt lång , eller hur ?
Tom vill bara vara lycklig .
Tom vet vad som pågår .
Tom skrattade åt Marys idé .
Tom lämnade vattnet på .
Tom lämnade kranen på .
Tom ljög för dig , eller hur ?
Tom ser upptagen ut , eller hur ?
Tom ser bra ut , eller hur ?
Tom gjorde sina föräldrar lyckliga .
Tom kan vara skadad eller död .
Tom nickade förstående .
Tom märkte Marys misstag .
Tom lade märke till skillnaden .
Tom pratar ofta med sig själv .
Tom öppnade kontorsdörren .
Tom lade sin hand på Marys .
Tom körde över någons hund .
Tom sa att han hade huvudvärk .
Tom sa att han var lycklig .
Tom sa att det här kunde hända .
Tom sa att du inte kunde komma .
Tom sa att du lät det hända .
Tom verkade riktigt förvirrad .
Tom verkar trivas här .
Tom verkar vara väldigt lycklig .
Tom borde inte vara härnere .
Tom borde inte ens vara här .
Tom öppnade långsamt dörren .
Tom stirrade på fotot på Mary .
Tom stirrade på dokumentet .
Tom studerade juridik på Harvard .
Tom lärde mig att köra bil .
Tom tror att det är omöjligt .
Tom trodde att du var full .
Tom sa att du tycker om hundar .
Tom sa att du var lycklig .
Tom tog ett foto på Mary .
Tom tog bussen till skolan .
Tom försökte öppna dörren .
Tom försökte öppna dörren .
Tom ville att jag skulle besöka honom .
Tom ville trösta Mary .
Tom var inte på Marys fest .
Tom var inte så säker själv .
Tom var själv inte så säker .
Tom gick ut genom bakdörren .
Tom skulle aldrig lämna Mary .
Tom är en mycket bra ingenjör .
det är snart Toms födelsedag .
Toms katt fick nio ungar .
Toms efternamn är Jackson .
Tom heter Jackson i efternamn .
Toms vänstra sko är borta .
Toms ben brändes svårt .
Toms lojalitet är beundransvärd .
Toms namn var på listan .
Tom är inte härifrån .
Tom är inte intresserad av matematik .
Toms föräldrar är lärare .
Toms svar överraskade Mary .
Toms berättelse förändras hela tiden .
det är Tom som är rädd .
Tom , jag måste prata med dig .
Tom , har du dina nycklar ?
Tom , titta vad du har gjort .
Tom , ring mig är du snäll .
Tom , du måste hjälpa mig .
vänta på din tur .
vi vet alla vad som kommer att hända .
vi gick också till templet .
vi bryr oss inte om vad han gör .
vi menar er inget illa .
vi har så mycket att diskutera .
vi måste handla .
vi måste göra det som är rätt .
vi måste fatta ett beslut .
vi måste börja nu direkt .
vi fattar beslut tillsammans .
vi behöver lite ljus härinne .
vi har bara tre alternativ .
vi har bara tre valmöjligheter .
det borde vi göra tillsammans .
det är bäst att vi gör som Tom säger .
det är bäst att vi inte åker fast .
vi kommer att behöva din hjälp .
vi kommer att bära gasmasker .
vi kommer att ta med mycket mat .
det tar vi hand om senare .
vi tar hand om dem senare .
vi tar hand om det här senare .
vi åker om en vecka idag .
vi åker om en vecka i dag .
vi måste jobba på det .
vi kommer aldrig att få veta vem han är .
vi kommer att ses igen .
vi ska tala om det där snart .
det ska vi tala om snart .
vi väntar tills det är mörkt .
vi är ute efter samma sak .
vi är nästan färdiga här .
vi är redan goda vänner .
det är vi som ställer frågorna .
vi är medvetna om problemet .
vi är bättre än de .
vi ska köpa mat åt dem .
vi kommer tillbaka imorgon .
vi kommer med dig , Tom .
vi följer med dig , Tom .
vi glömmer en sak .
vi tänker ge dig huset .
vi åker tillbaka till Boston .
vi ska gå på Toms fest .
vi kommer att vara tillsammans .
vi ska ändra på det .
vi ska göra vårt bästa .
vi ska hitta ett botemedel .
vi ska slutföra det här .
vi ska gifta oss .
vi ska spela ett spel .
vi ska leka en lek .
vi ska gå och spela tennis .
vi ska skydda dig .
vi ska äta biff ikväll .
vi är på väg tillbaka till stan .
vi är i samma bransch .
vi söker en advokat .
vi gör ett stort misstag .
vi gör inte det här igen .
vi är inte ens gifta ännu .
vi är inte härifrån .
vi går inte tillbaka dit .
vi tänker inte göra det .
vi tänker inte sälja den .
vi kommer inte att sälja den .
vi är inte här för att ha roligt .
vi tänker inte lämna dig här .
vi är inte tillsammans längre .
vi försöker spara pengar .
vi måste ta risken .
vi har väldigt lite tid på oss .
vi har aldrig gjort det förut .
vi har bara tre timmar på oss .
vi har sett vad Tom kan göra .
vi har sett vad du kan göra .
vi har sålt alla biljetter .
nå , vad är du bra på ?
det Tom såg överraskade honom .
vad gör vi här ute ?
vad trodde Tom att du gjorde ?
vad sa de att hade hänt ?
vad gjorde du i går kväll ?
vad matade du hunden med ?
vad vet du om honom ?
vad tror du att hände ?
vad vill du ska hända ?
vilken effekt kommer det att ha ?
vad hände egentligen här ?
vad var det som hände här egentligen ?
vad har hänt med din hand ?
vad är det du tror att jag gjorde ?
vad är ditt modersmål ?
vad gjorde du egentligen ?
vad skulle du vanligtvis göra ?
vad tänker du på ?
vilken är din favoritfilm ?
när kan jag komma härifrån ?
när byggdes det här templet ?
Varifrån fick du äggen ?
var bor din morbror ?
var bor din farbror ?
var finns det en telefon ?
var jobbade Tom då ?
vart skulle du vilja åka ?
vilken våning bor du på ?
vem vill du prata med ?
vem är det som äger pistolen ?
vem mer kom till festen ?
vem gav dig det här dokumentet ?
vem uppfanns telefonen av ?
vem sa att jag stal pengarna ?
vem körde likbilen ?
vem fattar besluten ?
varför ser du så ledsen ut ?
varför är du så trött idag ?
varför gjorde Tom så som han gjorde ?
varför tog du med Tom hit ?
varför tog ni med Tom hit ?
varför kom du tillbaka hit ?
varför behöver du de här pengarna ?
varför behöver du dessa pengar ?
varför vill du sälja den ?
varför vill du sälja det ?
varför vill ni sälja den ?
varför vill ni sälja det ?
varför går inte människor i ide ?
ska vi inte gå ut och äta ?
varför har du inte klänning på dig ?
ta på dig en klänning då .
varför beter sig Tom på det här sättet ?
kvinnor förtjänar jämställdhet .
andra världskriget tog slut 1945 .
vill du att jag ska köra ?
skulle du hellre stanna här ?
skulle ni hellre stanna här ?
Skriv med en kulspetspenna .
du klagar alltid .
du kan lämna rummet nu .
du visste att det här kunde hända .
du vet att det här är annorlunda .
du ser ut som Harry Potter .
du borde gå till tandläkaren .
du sa att Tom var annorlunda .
du sa att du var läkare .
du borde ha slutat tidigare .
du borde inte vara tillbaka här .
du borde inte vara här bak .
du borde inte ens vara här .
du är allt bra dum .
du börjar tråka ut mig .
du måste följa med mig .
ni måste följa med mig .
din fråga är ologisk .
din skjorta är inte instoppad .
ett glas rödvin , tack .
en tredjedel är mindre än en halva .
är du alldeles säker ?
är du för eller mot det här ?
är du ledig i eftermiddag ?
är du redo för Halloween ?
är du säker på att det är säkert ?
är ni säkra på att det är säkert ?
försöker du stöta på mig ?
Peking är större än Rom .
Beijing är större än Rom .
Småkryp attraheras av ljus .
men varför är det hela så hemligt ?
förresten , hur gammal är du ?
förresten , hur gamla är ni ?
kan jag tala med dig en sekund ?
kan vi åka nu ?
kan vi prata franska istället ?
skulle du kunna rita en karta åt mig ?
skulle du kunna ta det här , tack ?
skulle du kunna ta den här , tack ?
visade han dig bilden ?
hade du en trevlig kväll ?
hade ni en trevlig kväll ?
gör det som gör dig lycklig .
vet ni vem Tom är ?
har du ett hus i Italien ?
har du några förslag ?
har du skor och strumpor ?
känner du till några grekiska myter ?
gillar du dem verkligen inte ?
lider du av sömnlöshet ?
tycker Tom om Earl Grey @-@ te ?
åker han buss till skolan ?
glöm inte era pass .
Franskan utvecklades från latin .
ut härifrån ! allihopa !
gå upp tidigt på morgonen .
Guld är tyngre än silver .
grekiska är svårt att lära sig .
har Tom berättat allt ?
har Tom berättat allt för dig ?
har du borstat tänderna ?
har du funderat på terapi ?
han kom tillbaks två dagar senare .
han kan inte ha tappat bort sina nycklar .
han dog i cancer förra året .
han är ett matematiskt geni .
han är alltid vänlig mot mig .
han gräver sin egen grav .
han åker om tre dagar .
han längtar efter stadsliv .
han längtar efter stadslivet .
han står på scenen .
han valde ut den bästa boken .
han sa att han inte visste .
han berättade sin livshistoria för mig .
han deltog i mötet .
hennes dröm är att besöka Paris .
hennes söner har åkt till Tokyo .
hans fel var avsiktligt .
hans stackars hund lever fortfarande .
hans fru dog i barnsäng .
hur lärde du känna henne ?
hur lärde du känna honom ?
vad tyckte du om den där filmen ?
hur firade du jul ?
hur firade ni jul ?
hur löser jag det här problemet ?
hur löser jag detta problem ?
hur långt ifrån havet är vi ?
hur länge har du känt Tom ?
hur länge har ni känt Tom ?
hur länge tänker du stanna här ?
jag håller med dig helt och hållet
jag spelar volleyboll nu .
jag kan inte göra det här utan dig .
jag kan inte göra det här utan er .
jag kan inte göra detta utan dig .
jag kan inte ens göra en omelett .
jag kan inte komma på texten .
jag kommer inte ihåg texten .
jag minns inte texten .
jag klandrar dig definitivt inte .
jag valde mellan två alternativ .
jag är säker på att jag hörde ett skrik .
jag vet inte ens vem han är .
jag har inte mycket pengar nu .
jag tycker inte om att se Tom ledsen .
jag åt snabbt upp min lunch .
jag antar att detta var oundvikligt .
jag hatar alla slags insekter .
jag har en bok om fiske .
jag har en fruktansvärd tandvärk .
jag har precis ätit färdig .
jag måste låna lite pengar .
jag måste tala om det för Tom .
jag har mycket låg självkänsla .
jag hörde någon skrika nyss .
jag hörde någon skrika alldeles nyss .
jag visste att vi skulle vinna .
jag vet exakt var Tom är .
jag vet exakt var Tom befinner sig .
jag vet att du saknar din familj .
jag lärde mig att läsa i skolan .
jag lånade ut en del pengar till min vän .
jag gillar ris mer än bröd .
jag gillar österrikisk musik .
jag tycker om österrikisk musik .
jag gör dig nervös , inte sant ?
jag gör er nervösa , inte sant ?
jag kanske är din enda vän .
jag behöver någon att prata med .
jag behöver förbättra min franska .
jag kunde aldrig hålla en hemlighet .
jag ser ofta på dokumentärer .
jag spelar tennis en timme om dagen .
jag såg en gammal vän .
jag såg någonting intressant .
jag trodde knappt mina ögon .
jag borde inte ha lagt mig i .
jag låg kvar i sängen hela morgonen .
jag tror jag vet vad det här är .
jag tänker på dig hela tiden .
jag tror att det är där Tom är .
jag tror att det är där Tom befinner sig .
jag tror att den här killen menar allvar .
jag trodde att Tom var i skolan .
jag trodde att Tom skulle komma .
jag trodde att Tom skulle dyka upp .
jag besöker honom varannan dag .
jag vill komma till hotellet .
jag vill åka tillbaka till Italien .
jag vill veta vad som är roligt .
jag vill veta vad som är så roligt .
jag vill veta vad det är som är roligt .
jag vill veta vad det är som är så roligt .
jag var kolugn .
jag var här när du kom in .
jag skulle precis gå hem .
jag skulle precis göra det .
jag tränar för att hålla mig i form .
jag skulle göra vad som helst för dig .
jag kommer tillbaka om tio minuter .
jag låter dig sköta snacket .
jag är sprickfärdig av nyfikenhet .
jag kommer att behöva din hjälp .
jag ska tänka på det .
jag får inte hjälpa dig .
jag måste kila till banken .
jag har aldrig sett en tjock vegan .
Island hörde till Danmark .
om du är trött , så gå och lägg dig .
om ni är trötta , så gå och lägg er .
tänker någon äta det där ?
är det någon som tänker äta det där ?
är det någon som kommer att äta det där ?
kommer någon att äta det där ?
är det nyttigt för dig att äta fisk ?
är det din nya flickvän ?
det var faktiskt inte så illa .
det regnade mycket den vintern .
det startade en kedjereaktion .
det var Tom som stack ned Mary .
det var ett väldigt spännande spel .
låt oss hoppas på bra resultat .
många tror att jag är tokig .
Mary hjälpte sin mor att laga mat .
Mary hjälpte sin mamma att laga mat .
skulle jag kunna få låna telefonen ?
pengar växer inte på träd .
de flesta tror att jag är galen .
de flesta tycker att jag är galen .
min franska är lite rostig .
min bror är äldre än jag .
min dotter tycker om äggulor .
Vänd aldrig ryggen mot Tom .
ingen bryr sig om vad du tycker .
ingen kommer att klandra dig .
ingen kommer att beskylla er .
det är tydligt att någon ljuger .
Åh nej ! mitt hus brinner !
vår värd erbjöd oss en drink .
det är roligt att måla påskägg .
att spela tennis är hans hobby .
var snäll och stäng av motorn .
var har bildats i såret .
Ställ bilen i garaget .
Rapporterna ska lämnas in kommande måndag .
ett flertal människor skadades .
hon blev polis .
hon köpte en kamera till sin son .
hon bestämde sig för att säga upp sig från sitt jobb .
hon gav mig inte sitt namn .
hon har inte många böcker .
hon gav honom en massa pengar .
hon har en papegoja som husdjur .
hon ser ung ut för sin ålder .
hon blir sen till maten .
hon kommer att betala för allting .
kort hår passar henne verkligen .
Vissa sjukdomar är obotliga .
Vissa tjejer lär sig aldrig .
säg vad problemet är .
tala om för mig vad problemet är .
tennis är min favoritsport .
tack för er gästfrihet .
tack för din gästfrihet .
det är det jag är så stolt över .
djuret dog av svält .
svaret missar poängen .
svaret hade markerats fel .
Pilen missade sitt mål .
den vackra kvinna är vänlig .
boken kostar fem dollar .
paret hade ett lyckligt liv .
paret levde ett lyckligt liv .
dödläget var ett faktum .
hunden hoppade över en stol .
hunden vill gå ut .
valet låg mycket nära .
valet var mycket jämnt .
det är varmt på ön hela året .
mannen satte eld på sig själv .
bilden är verklighetstrogen .
priset är inte rimligt .
det har blivit mulet .
Ränderna var vågräta .
Förhandlingarna borde börja snart .
teven fungerar inte .
deras skepp ligger fortfarande i hamn .
det finns mjölk i kylen .
det fanns inga tecken på liv .
det finns inte mycket mer att tillägga .
det finns rum för diskussion .
det finns utrymme för diskussion .
det lämnas utrymme för diskussion .
de vill inte att du ska veta .
de gick mot porten .
de gick och fiskade i går .
de stod på rad .
denna bok verkar intressant .
jag förstår mig inte på det här .
den här flaggan är mycket vacker .
det här är Toms favoritbok .
det här är en turkisk tradition .
detta kommer att ta år .
det här kommer att ta år .
detta kommer att ta åratal .
det här kommer att ta åratal .
det här är verkligen inte rätt tillfälle .
det är här som Tom brukar hänga .
det här är Tom brukar hänga .
Tom blev nästan påkörd av en bil .
Tom och Mary adopterade en flicka .
det går bra för Tom och Mary .
Tom frågade om han var inbjuden .
Tom frågade om han var bjuden .
Tom gjorde det mot sin vilja .
Tom gjorde det mot hans vilja .
Tom tycker inte om grapefrukt .
Tom kom näst sist .
Tom hittade pengarna som saknades .
Tom hittade de försvunna pengarna .
Tom hittade pengarna som var borta .
Tom fick Mary att laga middag .
Tom fick schampo i ögonen .
Tom hade massor av frågor .
Tom har för mycket arbete att göra .
Tom är fullkomligt skräckslagen .
Tom är rädd för Marys hund .
Tom är alltid full av idéer .
Tom är en illegal invandrare .
Tom är väldigt hemlighetsfull .
Tom är duktig i skolan .
Tom är gift med en lärare .
Tom syns inte till någonstans .
Tom är ganska oansvarig .
Tom är smartare än Mary .
Tom är fortfarande rädd för Mary .
Tom är inte lika gammal som Mary .
Tom vet Marys hunds namn .
Tom vet vad Marys hund heter .
Tom lämnade hatten i bilen .
Tom gillar att läsa tidningar .
Tom tycker om te med kanel i .
Tom älskar mig , och jag älskar honom .
Tom öppnade skjutdörren .
Tom räfsade upp alla löv .
Tom insåg att Mary hade rätt .
Tom fyllde på sin kaffemugg .
Tom verkade vara väldigt imponerad .
Tom verkar vara intelligent .
Tom skickade Mary en inbjudan .
Tom skakade hand med alla .
Tom bodde i ett billigt hotell .
Tom stannade i ett billigt hotell .
Tom försökte begå självmord .
Tom går vanligtvis till skolan .
Tom ville gå på en promenad .
Tom ville ta en promenad .
Tom blev attackerad av en haj .
Tom attackerades av en haj .
Tom var helt hjälplös .
Tom var inte det minsta intresserad .
Tom är här vilken sekund som helst .
Tom arbetar från nio till fem .
Tom jobbar från nio till fem .
Tom har en tendens till att överdriva saker och ting .
två gånger sju är fjorton .
Vattenkraft roterar hjulet .
vi ska ha barn .
vi gick till konserten båda två .
vi kan ändra på oss om vi vill .
till slut gjorde vi upp en affär .
vi hade inget bättre för oss .
vi måste städa vårt klassrum .
vi studerade franska i skolan .
vi tycker att ni borde komma in .
vi kommer alltid att vara tillsammans .
vi skulle vilja ha en flaska rosé .
det Tom gjorde var otroligt .
vad tänker du på ?
vad gjorde du förra söndagen ?
vad föreslår du istället ?
vad tror du att det här är ?
vad vill du berätta för oss ?
vad gör vi om Tom inte klarar av det ?
vad händer om mina föräldrar får reda på det ?
hur är den nya ledaren ?
vad i hela världen står på ?
vilket skepp kom Tom med ?
vad är ditt modersmål ?
vad är ert modersmål ?
när flyttade du till Berlin ?
var är dina barn nu ?
var är era barn nu ?
var går Tom i skolan ?
var i Turkiet bor du ?
vilken webbläsare använder du ?
vem vill du prata med ?
vem vill ni prata med ?
vem vill du tala med ?
vem vill ni tala med ?
Vilka vill du tala med ?
Vilka vill du prata med ?
Vilka vill ni prata med ?
vem mer var på Toms fest ?
varför lyssnade du inte på mig ?
varför lyssnade ni inte på mig ?
skulle du vilja ha en till öl ?
skulle ni vilja ha en till öl ?
skulle du vilja ha en öl till ?
skulle ni vilja ha en öl till ?
du kan avbryta sökandet .
du får inte komma för sent den här gången .
du kan inte komma för sent den här gången .
ni kan inte komma för sent den här gången .
du får inte komma för sent denna gång .
ni får inte komma för sent denna gång .
du kan inte stanna här i natt .
du kan inte stanna här i kväll .
du måste inte göra det nu med en gång .
ni måste inte göra det nu med en gång .
det måste inte göras nu med en gång .
du måste städa ditt rum .
du måste vara jättehungrig nu .
du måste vara mer försiktig .
du behöver bara be om det .
ni behöver bara be om det .
ni behöver bara be om den .
du behöver bara be om den .
det borde du veta vid det här laget .
det var det här du ville , eller hur ?
din fråga har inget svar .
er fråga har inget svar .
&quot; hon gillar musik &quot; . &quot; det gör jag med &quot; .
faktiskt så är jag inte särskilt säker .
alla mina bröder har arbeten .
kan jag få komma med ett förslag ?
barn tycker om att klättra i träd .
Välj tre böcker på måfå .
kom tillbaka så snart du kan .
kan jag få ett glas vin ?
Brottslingar borde straffas .
Danzig är ett heavy metalband .
visade hon dig bilden ?
vet vi med säkerhet att det är Tom ?
vill du ha någonting att äta ?
vill du ha något att äta ?
vill du ha nåt att äta ?
vill du ha de där pralinerna ?
vill du se ditt rum ?
titta inte ut genom fönstret .
vill du inte simma idag ?
vill ni inte simma idag ?
Guds vägar äro outgrundliga .
har brevbäraren redan kommit ?
har du någonsin kysst en kvinna ?
har du någonsin sett den här flaggan ?
har du lärt dig din läxa ?
han högg ned det där körsbärsträdet .
han tyckte inte att det var kul .
han steg upp tidigare än han brukar .
han steg upp tidigare än vanligt .
han steg upp tidigare än normalt .
han hade massor att göra .
han skyndade sig tillbaka från England .
han är alltid snäll mot djur .
han kommer jämt för sent till skolan .
han kommer alltid för sent till skolan .
han klagar jämt och ständigt .
han är min bror , inte min far .
han kysste mig på pannan .
han lämnade allting åt slumpen .
han lade boken på hyllan .
han sa att han inte vet .
han stannade där hela tiden .
han kastade ut mig ur huset .
han opererades i går .
hennes syster bor i Skottland .
hans nya film är sevärd .
hur kan jag lösa det här problemet ?
hur kan jag lösa detta problem ?
hur länge har det snöat ?
hur länge har de varit här ?
hur mycket tjänar Tom ?
jag beundrar honom för hans mod .
jag ser alltid på dokumentärer .
jag tittar alltid på dokumentärer .
jag försöker att lära mig engelska .
jag försöker lära mig engelska .
jag bad henne att vänta ett slag .
jag tror att hon är ärlig .
jag kan inte låta det hända .
jag kunde inte fortsätta ljuga för Tom .
jag kräver en ursäkt från Tom .
jag drack inte te igår .
jag hjälpte mer än gärna till .
jag ville egentligen inte hjälpa till .
jag ville inte att det här skulle hända .
jag känner inte för att äta just nu .
jag vet inte vad klockan är .
jag känner inte riktigt för att dansa .
jag rekommenderar inte att göra det där .
jag tror inte att det här är tillräckligt .
jag förstår det inte heller .
jag vill inte gå till skolan .
jag hade en hamster som hette Cookie .
jag hade en hamster vid namn Cookie .
jag avskyr att se djur lida .
jag har en svår smärta i ryggen .
jag måste skriva några brev .
jag hoppas att ingen såg mig dansa .
jag hoppas att ni hade en trevlig resa .
jag vet att jag borde ha gjort så .
jag vet att Tom inte är lycklig där .
jag vet när din födelsedag är .
jag lärde mig att skriva i skolan .
jag lämnade en lapp under dörren .
jag vet bara vad Tom berättade för mig .
jag talar bara lite franska .
jag kan bara lite franska .
jag ville bara prata med Tom .
jag minns att jag mötte drottningen .
jag vinkade av honom vid flygplatsen .
jag tittar sällan på dokumentärer .
jag tycker att Tom borde varnas .
jag tycker att Tom är envis .
jag tycker att det är en dum idé .
jag tror att vi har tillräckligt med pengar .
jag trodde att Tom skulle komma ihåg .
jag trodde att Tom skulle minnas .
jag trodde att Tom skulle säga det .
jag tänkte att det var värt ett försök .
jag trodde du hatade rödvin .
jag trodde att du var annorlunda .
jag trodde att ni var annorlunda .
jag vill dricka en kopp te .
jag vill att du läser den här boken .
jag längtade efter en cigarett .
jag höll på att titta på en dokumentär .
jag såg en gammal film på tv .
jag åkte flygplan till Kyushu .
jag åkte till Kyushu med flygplan .
jag önskar att jag var lika lång som Tom .
jag undrar vem som namngav detta skepp .
jag skulle göra vad som helst för kärleken .
jag skulle vilja studera arabiska .
jag skulle vilja gå på bio .
jag skulle vilja ha två kilo äpplen .
jag skulle helst inte vilja sjunga idag .
jag sjunger helst inte i dag .
jag börjar ana ugglor i mossen .
jag går inte på mötet .
jag tänker inte gå på mötet .
jag är kapten över detta skepp .
jag har gjort allt jag kan för dig .
jag har lagat radion åt honom .
jag har aldrig varit i Argentina .
är det moraliskt fel att äta kött ?
det kvittar mig lika .
det är ett väldigt farligt system .
det är deras problem , inte vårt .
Japan är ett vackert land .
att lära sig koreanska är svårt .
vi sticker imorgon
Mary stängde tyst dörren .
får jag låna din ordbok ?
män vet inget om kvinnor .
de flesta barn älskar glass .
de flesta människor är högerhänta .
min ordbok är mycket användbar .
min farfar tycker om att promenera .
min morfar tycker om att promenera .
min farfar gillar att promenera .
min morfar gillar att promenera .
det gör ont i knät när jag böjer på det .
inget mer , tack . jag är mätt .
inga av de här äggen är färska .
inget är omöjligt för Gud .
nu har de tre barn .
ett språk är aldrig nog .
ett språk är aldrig tillräckligt .
våra mammor är starka kvinnor .
Känn dig som hemma .
Känn er som hemma .
var snäll och spika igen fönstren .
rödvin passar bra till kött .
hon började prata med hunden .
hon har en stuga vid havet .
hon har marginaliserat sig själv .
hon har platinablont hår .
hon är mer vis än smart .
hon var frånvarande på grund av en förkylning .
hon var på väg att svimma .
hon var svimfärdig .
hon var nära att svimma .
hon var på vippen att svimma .
efter söndag kommer måndag .
berätta för Tom vad du vill göra .
det låter som en bra överenskommelse .
det låter som en bra idé .
det är faktiskt en bra poäng .
det är inte riktigt mitt problem .
det är sant , jag lovar .
det är det vi väntar på .
det är det som vi väntar på .
pojken tittade in i rummet .
pojken gjorde sig lustig över flickan .
bilen körde in i ett skyddsräcke .
bilen satt fast i leran .
Bottenvåningen var översvämmad .
marknaden öppnar klockan nio på morgonen .
planet flög över Fuji .
det ligger en bok på bordet .
det finns ett piano i rummet .
det står ett piano i rummet .
det finns blott ett alternativ .
det finns ingen ost kvar .
det fanns ingenting i lådan .
det fanns inte en själ i sikte .
det är ingen stor skillnad .
de fångade rävar med fällor .
de bildade en ny regering .
de har ingen annanstans att ta vägen .
de skyndade sig ut ur rummet .
de talar spanska i Mexiko .
den här ölen är inte tillräckligt kall .
den här ölen är inte kall nog .
det här är Toms idé , eller hur ?
det är ett otroligt resultat .
det här är mycket viktigt för oss .
det är här vi båda hör hemma .
den här metoden är långsam men säker .
den här klockan var ett riktigt fynd .
den här jakten är väldigt dyr .
den här yachten är väldigt dyr .
denna lustjakt är väldigt dyr .
Tom har nästan aldrig på sig hatt .
Tom bär nästan aldrig hatt .
Tom bad mig klippa hans hår .
Tom åt en handfull russin .
Tom undvek militärtjänstgöring .
Tom hade knappt tillräckligt att äta .
Tom började bli nedstämd .
Tom kan inte bestämma sig för vad han ska köpa .
Tom kunde inte kontrollera sig själv .
Tom gjorde det för tre veckor sedan .
Tom gillade inte sin macka .
Tom vet inte att du är här .
Tom har inte ofta på sig hatt .
Tom bär inte ofta hatt .
Tom gillar inte riktigt Mary .
Tom tycker inte riktigt om Mary .
Tom gav Mary lite choklad .
Tom gav mig kikaren .
Tom har bevisat att det fungerar .
Tom har bevisat att den fungerar .
Tom har bevisat att det går .
Tom är professor i kemi .
Tom är en person som man kan lita på .
Tom ligger på en stor sten .
Tom jobbar på bilverkstan .
Tom jobbar på bilverkstaden .
Tom lämnade tv:n på hela natten .
Tom drog en suck av lättnad .
Tom tappade bort sin franska lärobok .
Tom tappade bort sin franska textbok .
Tom gillar verkligen inte Mary .
Tom tycker verkligen inte om Mary .
Tom rev upp kuvertet .
Tom sa att han inte äter kött .
Tom sade att han inte äter kött .
Tom dukade bordet för kvällsmaten .
Tom dukade bordet för middag .
Tom dukade för middag .
Tom sköt sig själv i knät .
Tom sover med strumporna på .
Tom dyker oftast upp i tid .
Tom var klädd helt i svart .
i morgon ska jag gå och shoppa .
vi tittade alla ut genom fönstret .
vi ska inte på semester .
vi kan inte lita på vad hon säger .
vi har inget annat val .
vi har inte tid för att debattera .
vi kände knappt dig på den tiden .
vi bor nära stationen .
vi måste gå tillbaka till skeppet .
vi föddes på samma dag .
vi går tillbaka till skeppet .
vi kommer att få det här gjort .
vi är väldigt tacksamma för det .
vi har talat om er .
det har varit en mycket svår vinter .
Tja , vad är det för fel med det ?
vilket företag jobbar du för ?
vilket företag jobbar du åt ?
vilket företag arbetar du för ?
vilket företag arbetar du åt ?
Vilka slutsatser kan vi dra ?
vilket är ditt favoritdjur ?
vilket skepp kommer du med ?
vad är problemet med det ?
vad gör den här stolen här ?
vilket är ditt favoritschampo ?
när behöver jag lämna tillbaka bilen ?
när borde jag lämna tillbaka bilen ?
var köpte du biljetten ?
var lärde du dig att skriva ?
Varifrån kommer pinjenötter ?
var finns närmaste toalett ?
vem vill ha lite varm choklad ?
varför ändrade du dig ?
varför är det ingen som hjälper Tom ?
du måste följa reglerna .
ni måste följa reglerna .
du sa att du var lycklig .
ni sa att ni var lyckliga .
du borde ha kommit med oss .
du borde slå upp det ordet .
du borde slå upp det ordet .
du berättar inte sanningen .
Bränt barn skyr elden .
faktiskt så hittade jag på det där .
Tillsätt naturell yoghurt och sojamjölk .
söker ni något ?
förresten , var bor du ?
var bor du , förresten ?
kan jag få lite varm choklad ?
kan du uttala de här orden ?
kan du visa mig en gång till ?
kan du inte stanna en stund till ?
stäng dörren när du går .
skulle ni kunna ge mig lite råd ?
trodde du verkligen det ?
kom du med första tåget ?
skrev du ned telefonnumret ?
titta inte ut genom fönstret .
känner du till någon bra restaurang ?
vet du hur man spelar schack ?
tycker du om chokladpudding ?
tror du att det kommer att regna idag ?
tror ni att det kommer att regna idag ?
vill du veta sanningen ?
var inte för sträng med dig själv .
bli inte så högfärdig .
torka byxorna på elementet .
ät din soppa medan den är varm .
det bor få människor på ön .
ge mig en till kopp kaffe .
ge mig något att skriva på .
ge mig tre kritor .
grekiska är inget enkelt språk .
grekiska är inget lätt språk .
Greker äter också mycket fisk .
har du packat klart än ?
har du pratat klart nu ?
han säger alltid samma sak .
han anlände tidigare än vanligt .
han kom fram tidigare än vanligt .
han kom hem senare än vanligt .
han trodde inte sina ögon .
han kunde inte gå längre .
han undersökte Amazonas regnskog .
han utforskade Amazonas regnskog .
han genomforskade Amazonas regnskog .
han fyllde glaset med vin .
han är alltid flitig som en myra .
han ber alltid om pengar .
han är en fullkomlig främling för mig .
han är stolt över att vara doktor .
han är stolt över att vara läkare .
han är längre än sin bror .
han lämnade boken på bordet .
han verkar inte ha vetat det .
han slog sig ner på en stol .
han sade till henne att han älskade henne .
hej , jag är Tom . vad heter du ?
hans tjänster uppskattades .
håll bollen med båda händerna .
vad sägs om en promenad på stranden ?
hur löste du problemet ?
hur säger man det på franska ?
hur länge har du varit utomlands ?
hur många böcker äger du ?
hur många månar har Mars ?
hur ska vi skydda oss själva ?
jag är en elev på den här skolan .
jag börjar komma ihåg det .
jag frågade honom vad han hette .
jag hör till basebollaget .
jag har inte råd att betala så mycket .
jag stannade inte där särskilt länge .
jag stannade inte särskilt länge där .
jag har ingenting att läsa .
jag har inga kläder att använda .
jag känner inga blinda .
jag vet inte om han är en doktor .
jag vet inte om han är en läkare .
jag vill inte prata om det .
jag tycker om att se på fotboll på tv .
ibland känner jag mig ledsen .
jag går till jobbet klockan sju .
jag fick ett brev från min vän .
jag fick en massa myggbett .
jag fick mig något att äta .
jag har många samtal att ringa .
jag har många beslut att fatta .
jag har varit i USA två gånger .
jag har levt här under en lång tid .
jag har mitt eget sovrum hemma .
jag hoppas att det ska vara bra imorgon .
jag hoppas att det är bra i morgon .
jag vet att hon har varit upptagen .
jag vet när någon ljuger för mig .
jag känner din bror väl .
jag lämnade mitt kreditkort hemma .
jag klarar av att försörja min familj .
jag har säkert ätit någonting konstigt .
jag skulle aldrig ha litat på Tom .
jag önskar bara att Tom vore här .
jag önskar bara att Tom kunde vara här .
jag spelade tennis hela dagen .
jag ångrar att jag åt ostronen .
jag borde sluta skjuta upp saker och ting .
jag klev på Toms hunds svans .
jag tar hand om min farfar .
jag tar hand om min morfar .
jag tror jag ska gå och lägga mig .
jag tycker att hon är en ärlig kvinna .
jag trodde inte att du kände Tom .
jag gick en konstkurs i fjol .
jag låg och vred mig hela natten .
jag tittar vanligtvis på dokumentärer .
jag vill vara en ärlig person .
jag vill vara mer självständig .
jag vill köpa en tjeckisk tröja .
jag vill äta kinesiska nudlar .
jag vill åka dit en gång till .
jag vill gå dit en gång till .
jag vill att du blundar .
jag var hemma nästan hela dagen .
jag tänkte precis på dig .
jag funderade på planen .
jag gick hem för att byta kläder .
jag hämtar dig efter jobbet .
jag önskar att jag hade ett eget rum .
jag önskar att jag hade ett rum för mig själv .
jag kommer inte att kunna betala för den .
jag kommer inte att kunna betala för det .
jag skulle gärna vilja åka till USA .
jag skulle vilja åka till USA .
jag ska äta lunch med Tom .
jag kommer att behöva lite hjälp med det här .
jag kommer att börja äta mindre kött .
jag kommer att skära ned på kött .
jag kommer att skära ner på kött .
jag kommer att sakna Tom så mycket .
jag är inte på humör just nu .
jag är inte så orolig för Tom .
jag är väldigt upptagen för tillfället .
jag har bett Tom att inte göra så .
jag har lärt Tom franska .
jag har aldrig ätit kinesisk mat .
jag har aldrig hört talas om den staden .
jag underskattade aldrig Tom .
jag har fortfarande mycket att lära .
var snäll och påminn mig om jag glömmer bort .
jag föddes i Boston faktiskt .
är det bra eller dåligt ?
är det vad du har i åtanke ?
har den här affären söndagsöppet ?
är din fru fortfarande i Amerika ?
det är faktiskt inte riktigt så enkelt .
den har för många nackdelar .
det är onormalt att äta så mycket .
det kommer att bli ganska kyligt .
det ligger bara några minuter bort .
det är oartigt att peka på folk .
det verkar som att jag har en lätt förkylning .
det var ett väldigt dumt beslut .
det var ett extremt grymt krig .
det var fantastiskt att jobba med Tom .
det var väldigt kallt den kvällen .
det är ungefär lika stort som ett ägg .
det är dags för mig att sova .
låt oss göra det någon annan gång .
låt oss att försöka lösa gåtan .
titta på mig när jag pratar med dig !
min engelska är inte alls bra .
min storebror är lärare .
varken Tom eller Mary kan simma .
ingen gjorde något annat än att dansa .
ingen får gå dit .
Oslo är Norges huvudstad .
lägg dina böcker i ditt skåp .
hon köpte en bok i affären .
hon har en del egna pengar .
hon är nästan sextio år gammal .
hon åkte till Kyoto , eller hur ?
någonting fruktansvärt har hänt .
var försiktig så att du inte blir förkyld .
tack för allt du gjort .
tack för informationen .
den där pojken talar som en vuxen .
sjön ser ut som ett hav .
det museet är värt att besöka .
det är faktiskt ganska smart .
det är faktiskt bra nyheter .
det är precis vad Tom vill .
det är mitt favorituttryck .
det är det som är kruxet .
det är därför jag är här , faktiskt .
Seine flyter genom Paris .
lådan är för tung för att lyftas .
Tränaren gav mig några råd .
experimentet var lyckat .
hotellet drivs av hans farbror .
hotellet drivs av hans morbror .
Förlusten var en besvikelse .
polisen hann ifatt honom .
den blyga pojken mumlade sitt namn .
tåget försenades av snön .
vattnet dränkte gatorna .
Kvinnorna nådde sitt mål .
där är en katt i köket .
det är en katt i köket .
det finns en katt i köket .
det finns yoghurt i kylen .
de här skorna är gjorda i Italien .
dessa skor är tillverkade i Italien .
de befarar att han kan vara död .
de har något gemensamt .
de gjorde en märklig upptäckt .
det sägs att man är vad man äter .
de tittade på teve .
de tittade på tv .
den här stolen är gjord av plast .
det här är ett mycket märkligt brev .
det här är en mycket märklig bokstav .
denna produkt är tillverkad i Italien .
den här produkten är tillverkad i Italien .
det här arbetet är inte på något sätt lätt .
Tokyo är huvudstad i Japan .
Tokyo är Japans huvudstad .
Tom har nästan alltid på sig en hatt .
Tom slog nästan ihjäl Mary .
Tom ringer mig nästan varje dag .
Tom kan tala flytande franska .
Tom kan tala franska flytande .
Tom kan prata flytande franska .
Tom kan prata franska flytande .
Tom kunde inte bestämma sig .
Tom ville inte tala med mig .
Tom ville inte prata med mig .
Tom har inte alltid hatt på sig .
Tom bär inte alltid hatt .
Tom hade ingen anledning att vara arg .
Tom har inget lokalsinne .
Tom har något i sin hand .
Tom har något i handen .
Tom har någonting i handen .
Tom är en duktig cricketspelare .
Tom ritar på ett skissblock .
Tom sa att han ville vara här .
Tom sade att han ville vara här .
Tom sa att han var oskyldig .
Tom tar yoga på stort allvar .
Tom tycker att det är tillräckligt bra .
Tom försökte förbättra stämningen .
Tom försökte höja stämningen .
Tom försökte rädda Marys liv .
Tom besökte Boston förra månaden .
Tom ville bli bonde .
Tom ville gå till stranden .
Tom ville äga en bokaffär .
Tom vill vara med på festen .
Tom vill bli brandman .
Tom var lite besviken .
Tom var en av de lyckligt lottade .
Tom svetsade ihop rören .
Tom skulle aldrig ha skadat dig .
Tom skulle aldrig ha skadat er .
Toms föräldrar kom hem tidigt .
Toms tal var riktigt roligt .
Toms tal var verkligen roligt .
tyvärr berättade ingen det för oss .
var det här någon annans idé ?
skulle det här vara roligt ?
vi kan inte fortsätta utan Tom .
vi åker och fiskar då och då .
vi sover vanligtvis i det här rummet .
vi röstade emot förslaget .
vi tänker flytta till Boston .
vi blir inte yngre .
vi blir inte yngre än så här .
vad äter du just nu ?
vad orsakade strömavbrottet ?
hur såg rånaren ut ?
varför lär du dig engelska ?
vad för fråga är det där ?
vad är klockan i Boston nu ?
det du fick lära dig är fel .
det ni fick lära er är fel .
vad är ditt intryck av Tom ?
var kom det där skeppet ifrån ?
var hörde du den historien ?
var är den japanska ambassaden ?
var ligger den japanska ambassaden ?
var är resten av pengarna ?
vilken buss går till flygplatsen ?
vem är brevet adresserat till ?
varför klev Tom in i den där bilen ?
varför skulle Tom vilja hjälpa oss ?
kan du hjälpa mig en minut ?
kvinnor behandlas annorlunda .
vill du ha lite mer nötkött ?
kan du släcka ljusen ?
kan du släcka stearinljusen ?
jag antar att du skulle kunna ha rätt .
du tycker inte ens om choklad .
du måste inte göra det nu .
du måste inte göra det där nu .
ni måste inte göra det där nu .
du behöver inte göra det där nu .
ni behöver inte göra det där nu .
du tillbringar för mycket tid ensam .
var på din vakt .
din födelsedag närmar sig .
en katt har en svans och fyra ben .
en hunds nos är väldigt känslig .
allt jag vill är att åka och fiska .
jobbar du fortfarande med Tom ?
arbetar du fortfarande med Tom ?
det tog inte lång tid innan månen kom fram .
Peking förändras så fort .
båda mina systrar är gifta .
får jag besvära om saltet ?
kan vi hyra en av de här båtarna ?
har du några minuter ?
kan du inte stanna lite längre ?
kan jag låna din gräsklippare ?
kan jag få titta på de där fotografierna igen ?
har alla gjort sin läxa ?
gjorde alla sin läxa ?
har alla gjort sina läxor ?
har du någon hostmedicin ?
har ni någon hostmedicin ?
tror du att ni kan få in mig ?
vill du äta lite middag ?
är det någon som vet vad som hände ?
köp inga fler presenter åt mig .
har du ingenting att göra ?
har inte du något att göra ?
har ni ingenting att göra ?
har inte ni något att göra ?
en evighet är en väldigt lång tid .
fyll i formuläret med kulspetspenna .
hälften av äpplena var ruttna .
han går alltid hemifrån klockan sju .
han löste korsordet med lätthet .
han har ett stort antal böcker .
han har ingen chans att återhämta sig .
han pressas alltid på pengar .
han är nöjd med sin nya bil .
han är världens rikaste man .
han föll aldrig för frestelsen .
han satte sig på bänken .
han kallades att vittna .
han låg och sov under trädet .
han gick och lade sig klockan tio som han brukar .
han är tillbaka om tio minuter .
hennes hår är långt och vackert .
hans frånvaro berodde på sjukdom .
hur dödade du kackerlackan ?
hur dödade ni kackerlackan ?
hur länge har du väntat ?
hur länge har du stått och väntat ?
hur många språk kan du ?
hur vill du ha ditt kaffe ?
jag är inte det minsta orolig .
jag kan inte besvara din fråga .
jag kan inte låta dem göra så här mot mig .
jag kan inte komma underfund med de här siffrorna .
jag fångade en vacker fjäril .
jag har inga böcker att läsa .
jag har inga nära vänner .
jag tror inte det är en bra idé .
jag vill inte vara din vän .
jag gav tillbaka hennes ordbok
jag har en hund som kan springa snabbt .
jag glömde mina bilnycklar .
jag har tre frågor till dig .
jag har tre frågor till er .
jag lade på och ringde henne igen .
jag bara älskar sådana saker .
ja ba älskar såna saker .
jag känner tjejen som spelar tennis .
jag gillar det , men jag älskar det inte .
jag hann dit i tid .
jag träffade henne på vägen till skolan .
jag behöver tänka på mina barn .
det trodde jag aldrig om dig .
jag öppnade asken . den var tom .
jag hämtade Tom på stationen .
jag plockade upp Tom på stationen .
jag antar att han kommer tillbaka snart .
jag trodde att vi var bästa vänner .
jag gick längs huvudgatan .
jag vill köpa en ordbehandlare .
jag vill ändra mitt utseende .
jag vill dricka något kallt .
jag åt några jordgubbar .
jag ska lära dig att spela schack .
jag önskar att jag kunde måla sådär .
jag skulle vilja ställa en fråga .
jag skulle vilja stanna en natt .
jag skulle vilja simma i den här floden .
jag går och köper lite choklad .
vi ses igen när vi är tillbaka på skeppet .
jag är på väg mot Boston nu .
jag är faktiskt här för att hjälpa dig .
jag försöker bara tjäna en slant .
jag är inte beredd att kompromissa .
jag är ledsen , men det är omöjligt .
jag väntar på dig på mitt rum .
jag har faktiskt aldrig varit full .
jag har läst ut boken .
jag har bott här hela mitt liv .
jag har sett en massa häftiga saker .
jag har sett en massa coola saker .
på våren blir dagarna längre .
är det vad du ville köpa ?
är det vad du ville säga ?
är det någon som kan svara ?
gör det vänstra ben fortfarande ont ?
det är tydligt att han är hemma .
det var ett misstag från deras sida .
det kommer antagligen att snöa i morgon .
Kiev är Ukranias huvudstad .
låt mig berätta för dig om fallet .
Mary köpte en blå slips till Tom .
Mary köpte Tom en blå slips .
Mary är intresserad av politik .
Memorera dikten till nästa vecka .
mina ansträngningar producerade inga resultat .
mina försök gav inga resultat .
min far lagade en trasig stol .
min favoritdans är tango .
ingen av oss talar franska .
Fetma är en nationell epidemi .
bara kärlek kan krossa ditt hjärta .
bara kärlek kan krossa hjärtat .
endast kärlek kan krossa ditt hjärta .
endast kärlek kan krossa hjärtat .
endast kärlek kan krossa ens hjärta .
Pandor bor i bambusnår .
Paris är Frankrikes huvudstad .
kanske var jag för hård mot Tom .
fysik är mitt favoritämne .
att spela tennis är jätteroligt .
sitt inte på den där bänken är du snäll .
var snäll och stäng av teven .
hallon är väldigt dyra .
Läs så många böcker som möjligt .
ska vi inleda mötet nu ?
ska vi påbörja mötet nu ?
ska vi sätta i gång med mötet nu ?
hon är väldigt rädd för ormar .
hon ser ut att vara full .
hon betalade för att gå på konserten .
hon tycker mycket om att skriva dikter .
hon var gråtfärdig .
hon hade hjärtformade örhängen .
hon är ungefär i min ålder .
borde jag köpa någonting till honom ?
spanska är hennes modersmål .
Sveriges befolkning växer .
simning är en form av träning .
det där låter inte särskilt artigt .
det var det jag tänkte säga .
båda svaren är felaktiga .
bägge svaren är felaktiga .
jorden är där vi alla bor .
sjukhuset öppnade förra månaden .
ungarna bytte basebollkort .
barnen bytte basebollkort .
barnen böt basebollkort .
Japans huvudgröda är ris .
Mötesrummet är på nedervåningen .
männen gick för att jaga lejon .
nästa dag var juldagen .
dagen därpå var juldagen .
följande dag var juldagen .
situationen var mycket komisk .
Förhandlingarna kommer att ta tre dagar .
Tigern rymde från djurparken .
Tornet kommer att rasa .
Tornet stod mitt ibland ruinerna .
det finns många floder i Indien .
det ligger en apelsin på bordet .
de är alla oskyldiga barn .
de röstade om motionen .
de kommer inte förrän imorgon .
de lider av malaria .
denna byggnad är gjord av sten .
den här stolen är väldigt bekväm .
den här dörren har svetsats fast .
den här dörren är fastsvetsad .
detta är en kamera tillverkad i Japan .
det här är en bild av min syster .
detta är ett väldigt komplext problem .
jag har svårt att tro på det .
det här är svårare än jag trodde .
det här är svårare än jag förväntade mig .
Locket hör till den där burken .
det här verkar för bra för att vara sant .
tre dagar senare var Tom död .
jag ska inte till skolan idag .
Tom och Mary avskyr varandra .
Tom köpte Mary lite choklad .
Tom köpte lite choklad till Mary .
Tom köpte lite choklad åt Mary .
Tom kom för att be oss om hjälp .
Tom kan skriva med båda händerna .
Tom spelar faktiskt inte mycket .
Tom dricker inte öl hemma .
Tom vet inte vad han ska beställa .
Tom har vanligtvis inte på sig hatt .
Tom är en främling i den här staden .
Tom rensar sin garderob .
Tom ska vara tillbaka idag på eftermiddagen .
Tom häller upp ett glas mjölk .
Tom är så mycket äldre än jag .
Tom ser alldeles skräckslagen ut .
Tom sade att mötet gick bra .
Tom säger att du är bra på tennis .
Tom borde ha varit här vid det här laget .
Tom trodde att ingen var hemma .
Tom vill prova ett nytt schampo .
Tom var alltid villig att hjälpa till .
Tom var alltid hjälpsam .
Tom var alltid tjänstvillig .
Tom hade tur som hittade sina nycklar .
tvätta händerna innan du äter .
vi kunde inte godta hans berättelse .
vi vill inte överbelasta Tom .
vi hade väldigt kul .
vi har ett väldigt allvarligt problem .
vi måste genast operera .
vi måste operera med det samma .
vi måste ta itu med det här problemet .
vi valde numret på måfå .
vi höll på att frysa ihjäl .
vi är så glada över att ha dig här .
vad gjorde Tom med pengarna ?
vad gjorde Tom av pengarna ?
vad gjorde du med den här boken ?
vad gjorde du av den där boken ?
vad fick du i julklapp ?
vad fick ni i julklapp ?
vad ska du med pengarna till ?
vad vill du ha i julklapp ?
vad vill ni ha i julklapp ?
vad innebär det att tänka stort ?
vad har du för stjärntecken ?
vad är ditt stjärntecken ?
vad kostar den här radion ?
vilken yogaställning är din favorit ?
när ska skeppet anlända ?
när ska skeppet komma fram ?
var ligger den australiska ambassaden ?
vem är kapten över det här skeppet ?
vem är kapten över detta skepp ?
vilken är din favoritsuperhjälte ?
vem är din favoritsuperhjälte ?
kan du förklara vad det här är ?
vill du ha lite mer sås ?
skulle du vilja bli min vän ?
kan du vara snäll och låsa dörren ?
kan ni vara snälla och låsa dörren ?
kan du låsa dörren är du snäll ?
kan ni låsa dörren är ni snälla ?
du missbrukar dina maktbefogenheter .
du behöver inte svara idag .
du gillar visst inte sashimi ?
du får bara prata engelska .
du måste ta buss nummer 12 .
du ser precis ut som din pappa .
du ser väldigt blek ut . mår du bra ?
du måste vänta på nästa buss .
du borde inte titta ner på honom .
du kommer att glömma bort mig förr eller senare .
ditt förslag är lite extremt .
&quot; vem är det ? &quot; &quot; det är din mor &quot; .
ett kuvert och ett frimärke , tack .
är du rädd för skräckfilmer ?
är du rädd för rysare ?
är du för eller emot planen ?
så vitt jag vet är han inte lat .
fåglar sjunger tidigt om morgonen .
kan vi prata med dig en sekund ?
det är bara två veckor till jul .
julen är bara två veckor bort .
blunda och sov .
gav du verkligen Tom pengar ?
hörde du vad jag sade till Tom ?
såg du blicken han gav mig ?
såg du gårdagens avsnitt ?
har du någon astmamedicin ?
vet du varför himlen är blå ?
tror du verkligen på spöken ?
tror du fortfarande att jag bluffar ?
vill du ha lite äggröra ?
påminner det här dig om någon ?
fråga inte , bara gör det .
ingenting ont som inte har något gott med sig .
efter regn kommer solsken .
fem gånger sju är trettiofem .
ge mig en dollar för boken .
är det någon här som har varit i Boston ?
har du ätit färdigt frukosten än ?
han erkände att han hade tagit mutor .
han frågade om jag gillar kinesisk mat .
han tror på det övernaturliga .
han kan tala franska och engelska .
han förklarade sin situation för mig .
han tvingade sig in i rummet .
han har faktiskt inte ätit kaviar .
han hatar att bli tillsagd att skynda sig .
han är en man att räkna med .
han är min bror , inte min far .
han sparkade honom medan han låg ner .
han såg ut som om han vore sjuk .
ofta kommer han inte till skolan .
han visade mig hennes foto i smyg .
han kommer att besöka oss en dag .
han är tre år äldre än henne .
hans svar är i princip ett nej .
vad sägs om att spela schack i kväll ?
hur tar jag mig till busshållplatsen ?
hur långt är det till nästa bensinstation ?
hur långt är det till nästa mack ?
hur länge måste jag stanna här ?
hur många språk talar du ?
hur mycket av det här är Toms fel ?
hur mycket av detta är Toms fel ?
hur ofta cyklar du ?
hur ofta tvättar du håret ?
jag är van vid att jobba hårt .
jag är van vid att arbeta hårt .
jag är rädd att jag åt något dåligt .
jag måste tyvärr gå nu .
jag är upptagen med maten för tillfället .
jag är inte det minsta förvånad .
jag gick faktiskt aldrig på högskola .
jag såg det faktiskt inte själv .
jag har inte tid att läsa böcker .
jag gör inte Mary lycklig längre .
jag ser inget problem med detta .
jag tror inte att jag kommer att åka till Boston .
jag vill inte öppna fönstret .
jag vill inte prata om henne .
jag ville bara ställa en fråga .
jag ville bara kolla min mail .
jag ville bara kolla min mejl .
jag visste att Tom inte skulle förlora .
jag tycker om mandlar , men inte jordnötter .
jag bor i Boston med min familj .
jag älskar varenda en av er .
om det bara var så enkelt .
jag önskar bara att det var så enkelt .
om det bara vore så enkelt .
jag spelade tennis med min bror .
jag vill verkligen veta sanningen .
jag ångrar att jag inte åkte dit .
jag ångrar att jag inte gick dit .
jag respekterar dig och dina åsikter .
jag såg Tom för mindre än en timme sen .
jag såg Tom för mindre än en timme sedan .
jag kan fortfarande inte riktigt tro det .
jag pluggade i kanske två timmar .
jag tycker att han är en skicklig person .
jag tror att de flesta skulle samtycka .
jag trodde att du skulle vara redo vid det här laget .
jag tog ut kakan ur ugnen .
jag förstår vad du säger .
jag förstår vad ni säger .
jag vill komma i kontakt med henne .
jag vill sova lite längre .
jag vill att du håller ditt löfte .
jag låg i koma i tre år .
jag var tvungen att göra någonting .
jag funderade på planen .
jag kompenserar för det nästa gång .
jag önskar att jag hade varit med henne då .
jag undrar vem som satte igång det där ryktet .
jag skulle vilja ha något att dricka .
jag skulle vilja gå och sova nu .
jag skulle aldrig ha gissat det .
det skulle jag aldrig ha gissat .
jag skulle vilja skicka dessa till Japan .
jag går hellre än att ta bussen .
jag kommer aldrig att glömma din vänlighet .
jag är faktiskt en väldigt bra förare .
jag har faktiskt kul ikväll .
jag ser inte fram emot det .
det är inte meningen att jag ska tala med dig .
jag är inte säker på om det här är rätt .
jag kommer antagligen att försöka igen .
jag är trött på att bli kallad lögnare .
jag är trött på dina dumma kommentarer .
jag ber om ursäkt för det sena svaret .
jag är nöjd med mitt köp .
jag har faktiskt aldrig spelat golf .
jag har alla de vänner som jag behöver .
jag har haft det jättetrevligt i Boston .
jag har precis kommit tillbaka från Sverige .
är lektionen redan slut ?
det har blivit märkbart kallare .
det blir inte svårt att göra .
det skulle inte göra någon skillnad .
det skulle inte spela någon roll .
det är jättekul att vara här i Boston .
det är onekligen den bästa metoden .
Klava överförenklar allting .
låt mig ta ditt blodtryck .
jag tycker inte att vi pratar om det något mer .
Mary är verkligen en riktigt söt tjej .
de flesta av våra anställda är unga .
min engelska är allt men inte bra .
min engelska är allt utom bra .
min cykel behöver lagas .
min hund följer efter mig överallt jag går .
min åsikt skiljer sig från din .
mitt sommarlov är över .
Herregud , jag tror inte det är sant .
i vår trädgård finns två körsbärsträd .
var snäll och stäng dörren efter dig .
hon översatte det ord för ord .
hon är frånvarande för att hon är sjuk .
hon är orolig över din säkerhet .
hon är orolig över er säkerhet .
håll käften , annars åker du ut .
jag tog en tupplur eftersom jag var trött .
någon har stulit alla mina pengar .
det är långt ifrån sommar än .
tio procent är mer än tillräckligt .
så där behandlar han mig jämt .
så där behandlar han mig alltid .
det där är poeten som jag träffade i Paris .
det är emot mina principer .
det går emot mina principer .
det är inte vad jag gick med på .
katten sover på soffan .
Kakorna är under bordet .
Branden var på första våningen .
flickan stirrade på dockan .
stegen var täckt med lera .
sjön är stor och vacker .
det sista tåget har redan farit .
ljudet kommer att väcka bebisen .
Gubben är blind på ena ögat .
den gamle mannen är blind på ena ögat .
rummet är i oklanderligt tillstånd .
skeppet har inte ens dockat än .
skeppet börjar sakta att röra på sig .
Tornet kan ses härifrån .
äntligen är vi två ensamma .
det är för mycket att göra .
det ligger en apelsin på bordet .
det var inga varningar överhuvudtaget .
det fanns lite dagg imorse .
det fanns ingen i rummet .
de här muffinsen är nybakade .
de är min farfars böcker .
de är min morfars böcker .
de fångade räven med en fälla .
de har inte kommit tillbaka hem än .
den här kameran är tillverkad i Tyskland .
det här är en bild på Toms fru .
detta är en bild på Toms fru .
det här är dåligt för miljön .
det här kommer att bli intressant .
det här blir intressant .
det här svärdet är i gott skick .
tiden är ute . lämna in era uppsatser .
Tom hittar alltid fel hos henne .
både Tom och Mary är från Kanada .
Tom och Mary hade kuddkrig .
Tom anlände i grevens tid .
Tom anlände trettio minuter sent .
Tom ville inte döda någon .
Tom försvann utan ett spår .
Tom vill inte verka svag .
Tom följer en strikt vegansk diet .
Tom har inga vänner att leka med .
Tom har inte några vänner att leka med .
Tom kommer också till festen .
Tom håller på att söka efter ett bättre jobb .
Tom väntar på dig där uppe .
Tom kysste Mary på pannan .
Tom behöver köpa en ny regnrock .
Tom visade Mary staden .
Tom visade Mary runt i staden .
Tom tackade Mary för hennes råd .
Tom ville lära sig att läsa .
Tom såg på hela tiden .
Tom tittade hela tiden .
Tom tittade på hela tiden .
Toms familj bor i Australien .
vi frågade honom vad han hette .
vi får inte många besökare här .
vi vill inte ha någonting från dig .
vi njöt av att simma i sjön .
vi fattar varje beslut tillsammans .
vi såg många skepp i hamnen .
vi såg barnet kliva på bussen .
vi såg barnet stiga på bussen .
vad gjorde du i skolan idag ?
vad gjorde du i skolan i dag ?
vad gör du för att få tiden att gå ?
vad gör du för att fördriva tiden ?
vad tror du hände här ?
vad tror ni hände här ?
vilken frukt tycker du bäst om ?
vad heter den här gatan ?
vilken är din favoritsvordom ?
när bröt andra världskriget ut ?
när klippte du dig senast ?
var hittade du den här bilden ?
var bor du just nu ?
var bor ni just nu ?
var ligger den australiska ambassaden ?
var var du när det hände ?
var var du när det inträffade ?
var finns den närmsta bensinstationen ?
var ligger närmsta bensinstation ?
var ligger närmaste bensinstation ?
vilken av de två är tyngst ?
Vilkendera är tyngre ?
varför låter du inte bara Tom hjälpa till ?
varför låter ni inte bara Tom hjälpa till ?
varför har ingen sagt någonting ?
vilda djur bor i regnskogen .
vill du ha fler kakor ?
vill du ha te eller något ?
skulle du vilja dansa med mig ?
skulle du vilja se på en film ?
du har ingen anledning att vara rädd .
du måste fånga djuret levande .
ni borde fråga honom om råd .
du använder verkligen mycket smör .
du döljer någonting för mig .
du är gammal nog att förstå .
din bror ber om hjälp .
ditt problem liknar mitt .
&quot; hur gammal är du ? &quot; &quot; jag är sexton år &quot; .
ett spädbarn sover i vaggan .
en tiger har rymt från zoot .
en tiger har rymt från djurparken .
det står ett äpple på bordet .
eftersom han ljög straffades han .
Berlin är Tysklands huvudstad .
förresten , vad är din adress ?
kan du hjälpa mig att laga min punktering ?
dinosaurier härskade en gång över världen .
Samtycker du med deras beslut ?
vet du vilken färg hon gillar ?
vet du vad hon tycker om för färg ?
vet du vad hon gillar för färg ?
vet du vilken dag det är i dag ?
vet du vem som har skrivit den här romanen ?
kör du ofta bil till arbetet ?
vill du gå någon annanstans ?
kasta inte stenar i älven .
har du någonsin ätit en bananpaj ?
han gråter alltid när han är full .
han bråkar jämt med sin fru .
han behandlar mig alltid som ett barn .
han har byggt sig ett nytt hus .
han räknade ut ljusets hastighet .
hon kom först i tävlingen .
han vill inte prata om det .
han somnade med radion på .
han har en bror och två systrar .
han driver alltid med mig .
han sparkade in bollen i mål .
han må vara rik , men han är snål .
han var nöjd med resultatet .
han var tillfreds med resultatet .
han var sjuk , så han kunde inte komma .
han var siste man att komma fram .
han väger mycket mera än förut .
han kommer att återvända till Japan en dag .
han torkade svetten från ansiktet .
han arbetar hårt året runt .
hennes far avled i förra veckan .
hans rum är alltid i ordning .
vad sägs om att sätta på en kopp te ?
hur många språk kan du tala ?
hur mycket är du redo att förlora ?
hur mycket är ni redo att förlora ?
hur mycket är du beredd att förlora ?
hur mycket är ni beredda att förlora ?
hur ofta tvättar du dina jeans ?
jag kan faktiskt inte svaret .
jag vet faktiskt inte svaret .
jag klarar inte av att se blod .
jag klarar inte av synen av blod .
jag klarar inte av sådan här musik .
jag kan inte stå ut med detta ljudet längre .
jag står inte ut med det här oljudet längre .
jag står inte ut med detta oljud längre .
jag sa inte att det inte var okej att äta .
jag klandrar dig inte för att du gör så .
jag bryr mig inte om vad de säger .
jag har ingen mobiltelefon längre .
jag vet inte hur man köper en biljett .
jag vet inte vad jag ska göra imorgon .
jag tycker inte om pizza , men det gör Tom .
jag tycker inte om att jobba på helger .
jag har inget emot att göra hushållssysslorna .
jag tror inte att jag ska gå på college .
jag förstår inte den här meningen .
jag jobbar vanligtvis inte på helger .
jag vill inte höra några ursäkter .
jag vill inte ta några risker .
jag äter frukost klockan åtta .
jag har fjärilar i magen .
jag har inte tid att göra mina läxor .
jag har seglat på Themsen en gång .
jag har inte så mycket pengar med mig .
jag vill bara att människor ska vara försiktiga .
jag vill bara att folk ska vara försiktiga .
jag vill bara ha någon att prata med .
jag visste att du skulle sansa dig .
jag visste att ni skulle sansa er .
jag visste att du skulle komma till besinning .
jag visste att ni skulle komma till besinning .
jag vet hur svårt det är att göra så .
jag bor intill leksaksaffären .
jag bodde i det här huset som barn .
jag gjorde ett dåligt misstag på provet .
jag behöver ställa er några frågor .
jag har bara femtio med rep .
jag lovar . jag kommer aldrig att göra det igen .
jag vill verkligen komma underfund med det här .
jag skulle bara ha gått rakt in .
jag trodde att jag sa åt dig att inte komma .
jag vill helst inte prata om det .
jag skulle vilja åka till Frankrike någon gång .
jag förlåter , men jag kommer aldrig att glömma .
jag ska av på nästa station .
jag är faktiskt ganska seriös .
jag fryser . kan jag stänga fönstret ?
jag letar efter en vän till mig .
jag är inte van vid att göra det .
jag kokar fortfarande råriset .
jag är säker på att jag rätt nummer .
jag är trött . jag går och lägger mig .
jag har aldrig mått så bra i hela mitt liv .
jag har aldrig mått så bra förut .
i skolan blev Tom ofta mobbad .
är det dyrare att äta nyttigt ?
kommer han hem klockan sex ?
är det säkert att simma i den här floden ?
kommer presidenten att avgå ?
finns det någon bank nära stationen ?
det tog nätt och jämnt en timme .
det var min tur att städa rummet .
det kommer att kosta minst fem dollar .
visst är det vackert väder ?
det har varit varmt de senaste dagarna .
det är enkelt att göra och det är billigt .
det är verkligen inte mödan värt .
Kenya blev självständigt 1963 .
låt oss glömma alltsammans , okej ?
malaria bärs av myggor .
han har kanske många flickvänner .
pengar är det sista han vill ha .
min bror och jag delade rummet .
min pappa är inte hemma just nu .
min pappa är starkare än din .
min pappa sopar garaget .
min vän är sjutton år .
min syster leker med en docka .
ingenting är så enkelt som det verkar .
inget är så enkelt som det verkar .
man måste dra gränsen någonstans .
en av dina knappar har lossnat .
Paris är en ganska dyr stad .
Skala äpplet innan du äter det .
var snäll och lämna mig i fred . jag är upptagen .
hon har tagit på sig alltför mycket arbete .
hon är inte så ung som hon ser ut .
hon spelade piano tillräckligt bra .
hon kvävde honom med en kudde .
Oljetillgångarna är inte oändliga .
berätta nånting om dig själv .
tack för att du hjälpte mig att reparera bilen .
tack för att du tog hand om min hund .
den där dunkudden ser dyr ut .
det var en liten missberäkning .
det där var väldigt hänsynsfullt av Tom .
det där var riktigt kul . gör det igen !
det där var riktigt roligt . gör det igen !
det var inte alls vad jag trodde .
romarna förföljde kristna .
katten sover på bordet .
katten på bordet sover .
Datorreparationen tog hela dagen .
Levnadskostnaderna har sjunkit .
det är väldigt lätt att ta sig till ön .
ljudet väckte mig från min sömn .
planet gjorde en perfekt landning .
skeppet var inte redo för strid .
den sjuka mannens liv är i fara .
Trafikljuset slog om till rött .
båda svaren är korrekta .
bägge svaren är korrekta .
de sårade kom med ambulans .
det är en papegoja i fågelburen .
det finns en annan möjlighet också .
det är något fel på dig .
det är de som vill gå .
efter filmen somnade de .
de förorsakade oss knappt några problem .
saker och ting började ordna sig för Tom .
detta barnet har växt upp normalt .
det här smakar typ som kyckling .
i dag mår jag mycket bättre .
Tom kände nästan inte igen Mary .
Tom frågade Mary om hon kunde hjälpa honom .
Tom förnekade att det var han som var tjuven .
Tom verkade inte överraskad alls .
Tom verkade inte det minsta överraskad .
Tom går inte till jobbet på söndagar .
Tom gillar inte Marys attityd .
Tom tycker inte om Marys attityd .
Tom vill inte prata med dig .
Tom har inte hatt på sig varje dag .
Tom förlät Mary på hennes dödsbädd .
Tom har betett sig väldigt konstigt .
Tom har aldrig sett Mary så arg .
Tom är faktiskt väldigt bra på att laga mat .
Tom sover , men Mary är vaken .
Tom står inför finansiella problem .
Tom är äldre än vad resten av oss är .
Tom är en av mina närmsta vänner .
Tom är väldigt sportintresserad .
Tom vet verkligen inte vad han ska göra .
Tom gick ner på knä för att se bättre .
Tom läser nästan inga böcker alls .
Tom sade att han gick dit för ett jobb
Tom borde inte ha ätit så mycket .
Tom tog av sig sin rock och sina handskar .
Tom har på sig hatt nästan varje dag .
Toms familj äter sällan tillsammans .
vi kan inte ge upp utan en kamp .
vi gjorde vad vi var tvungna att göra för att överleva .
vi gjorde vad vi måste för att överleva .
vi vill inte vänta längre .
vi spelade schack och hade det trevligt .
vi måste respektera lokala seder .
vi måste prata med er om Tom .
vi måste prata med dig om Tom .
vi måste tala med er om Tom .
vi måste tala med dig om Tom .
vi satt mitt i rummet .
vi blev tillsagda att stanna på skeppet .
vi är tacksamma för er vänlighet .
vi är tacksamma för din vänlighet .
vi har gått runt hela sjön .
vad gjorde du i helgen ?
vilket tåg tänker du ta ?
vad är lufttemperaturen idag ?
vilket nagellack är din favorit ?
vilket är ditt favoritnagellack ?
varför hälsar Tom aldrig på oss längre ?
varför skulle någon vilja göra det ?
ord kan inte beskriva skönheten .
du får prata hur mycket du vill .
du måste alltid göra det rätta .
ni måste alltid göra det rätta .
ni ska alltid göra det rätta .
du har faktiskt rätt i det .
du är i bättre form än jag .
du har bättre kondition än jag .
ett DNA @-@ test visade att han var oskyldig .
med lite språkkunskaper kommer man långt .
en ekorre gömde sig bland grenarna .
Anpassning är nyckeln till överlevnad .
alla eleverna kommer från USA .
är du nöjd med resultatet ?
är du säker på att det här är Toms kontor ?
är du säker på att detta är Toms kontor ?
klarar du dig ensam i helgen ?
kan du hämta mig på stationen ?
kan ni hämta mig på stationen ?
kan du berätta vilken storlek den här är .
Kriminalitet lönar sig inte i längden .
Kriminalitet lönar sig inte i det långa loppet .
Kriminalitet lönar sig inte på lång sikt .
hade du roligt i helgen ?
går det bra att jag sänker volymen på teven ?
äter du ofta fisk till middag ?
gillar du verkligen inte de där killarna ?
vill du se det här programmet ?
tycker din flickvän om blommor ?
förvänta dig inte att alla ska tycka om dig .
förvänta dig inte att alla ska gilla dig .
glöm inte vad jag nyss sa till dig .
glöm inte vad jag nyss sade till dig .
glöm inte vad jag nyss sa till er .
glöm inte vad jag nyss sade till er .
glöm inte vad jag sade till er nyss .
glöm inte vad jag sa till er nyss .
glöm inte vad jag sa till dig nyss .
glöm inte vad jag sade till dig nyss .
kasta ingenting på marken .
alla vill sitta bredvid henne .
som tur är var vädret bra .
Lyckligtvis var vädret bra .
som tur var , var vädret bra .
Gud skapade jorden på sex dagar .
Gud skapade världen på sex dagar .
Greta Garbo var en svensk skådespelare .
har du någonsin ätit japansk mat ?
har du inte diskat än ?
han bedrog sina vänner för pengar .
han skar upp köttet och vägde det .
han beskrev flygresan i detalj .
han talade inte såvida han inte blivit tilltalad .
han drack direkt ur flaskan .
han tjänar tre gånger så mycket som jag .
han har ett stort hus och två bilar .
han har det bättre än någonsin .
han gillar matematik , men det gör inte jag .
han letade efter dem i fem timmar .
han satt där med sina ögon stängda .
han visade mig hennes bild i smyg .
han borde ha varit färdigt nu .
han var rädd att du skulle skjuta honom .
han kommer kunna gå upp och gå om ungefär en vecka .
hur ska Tom ta sig ur det här ?
jag tycker inte om honom , men jag gillar henne .
jag vet inte vad det här ordet betyder .
jag vet inte vad jag ska öppna den med .
jag vet inte vad jag ska öppna det med .
jag gillar inte att bli driven med .
jag minns inte vad han heter .
jag vill inte träffa någon i dag .
jag gav dem ett tusen yen var .
jag har en vän vars namn är Tom .
jag har en vän som heter Tom .
jag har aldrig ätit mango förut .
jag har inte försökt göra det på det sättet .
jag hörde Tom sjunga i duschen .
jag vet att det där inte är Toms underskrift .
jag tycker om att läsa innan jag går och lägger mig .
jag tycker bättre om vitt vin än rött .
jag uppskattar verkligen din hjälp .
jag uppskattar verkligen din vänlighet .
jag minns allt du säger till mig .
jag tror att jag måste skaffa nya glasögon .
jag tror det är dags för mig att dra .
jag trodde att Tom skulle vara på baren .
jag trodde aldrig att Tom skulle hålla käften .
jag tog mig friheten att ringa henne .
jag försöker att aldrig äta efter klockan åtta .
jag uppskattar vår vänskap mycket .
jag vill ha en massage . jag behöver slappna av .
jag var försenad på grund av trafiken .
jag var tillsammans med vänner hela förra natten .
jag åkte till flygplatsen för att träffa honom .
jag åkte till flygplatsen för att möta upp honom .
jag önskar att Tom var här med mig idag .
jag önskar att Tom var här med oss idag .
jag undrar vems sax det här är .
jag skulle vilja ringa ett samtal .
jag skulle vilja sova lite längre .
jag tar en kopp kaffe , tack .
jag är egentligen en universitetslärare .
jag börjar tappa tålamodet .
jag ska delta i en demonstration .
jag ska gå med i en demonstration .
jag ska träffa en kompis efter skolan .
det är inte meningen att jag ska göra detta .
jag är världens lyckligaste man .
det var jag som lärde Tom franska .
jag har aldrig hört den är låten innan .
om jag var rik så skulle jag åka utomlands .
om jag vore rik , skulle jag åka utomlands .
säg till om du är trött .
säg till om ni är trötta .
säg till om du blir trött .
säg till om ni blir trötta .
är det tufft att jobba på McDonald &apos; s ?
är det något fel på dina ögon ?
är din lägenhet väl underhållen ?
det har aldrig snöat på ön .
hon kommer förmodligen .
det är verkligen inte mödan värt .
det var en obeskrivlig situation .
det är normalt att vara lite rädd .
det är inte blod . det är tomatsås .
håll ett öga på min väska en stund .
håll ett öga på min väska ett slag .
Sömnbrist är inte bra för kroppen .
låt oss klä granen .
vi klär granen .
vi klär julgranen .
låt oss klä julgranen .
vi sätter julgranen här .
vi ställer julgranen här .
Mary satte några blommor i vasen .
min familj är väldigt viktig för mig .
ingen medicin kan bota denna sjukdom .
ingen medicin kan bota den här sjukdomen .
inga stjärnor syntes på himlen .
vår fotbollsmatch kommer att skjutas upp .
snälla be Tom att säga sanningen .
hon vill inte prata om det .
hon har känt honom länge .
hon har många vänner i Hong Kong .
hon skadades i en bilolycka .
hon bar en vacker klänning .
några barn leker i parken .
Vissa kvinnor rakar inte benen .
Vissa kvinnor rakar inte sina ben .
Somliga kvinnor rakar inte benen .
Somliga kvinnor rakar inte sina ben .
någon stal mitt körkort .
ibland förstår jag mig inte på honom .
ibland förstår jag inte honom .
ibland förstår jag honom inte .
det är lättare att lyfta än att landa .
tio är tio procent av etthundra .
1,6 mil är inte en kort sträcka .
tack så mycket för att ni bjöd in mig .
tack så mycket för att du bjöd in mig .
det skulle inte spela någon roll .
det där är anledningen varför han blev arg .
det är anledningen till att han blev arg .
det är orsaken till varför vi skilde oss .
djuret gav ifrån sig ett gnällande ljud .
kommittén sammanträder två gånger om månaden .
kommittén sammanträder två gånger i månaden .
kommittén sammanträder två gånger per månad .
jorden är mindre än solen .
familjen åt sin middag vid tolv .
gruppen springer på stranden .
Parkeringsplatsen är gratis .
Upprorsmännen saboterade järnvägen .
rebellerna saboterade järnvägen .
rummet kommer att målas imorgon .
Våldet varade i två veckor .
det finns femtio stater i Amerika .
Amerika har femtio stater .
det ligger affärer längs gatan .
det finns en tv i rummet .
det var ingen där förutom jag .
det fanns ingen där förutom jag .
det finns inte en chans att jag går in dit .
de lade ut mattan på golvet .
det här kaffet smakar diskvatten .
det här är en bild på Toms familj .
detta är en bild på Toms familj .
det här är brevet från min vän .
den här medicinen kommer att bota din förkylning .
Tom och jag , vi båda saknar dig väldigt mycket .
Tom och Mary väntade inte på John .
Tom frågade Mary varför hon var så arg .
Tom verkar inte komma åt sina data .
Tom verkar inte komma åt sin data .
Tom kom inte hem förrän vid midnatt .
Tom glömde att ställa väckarklockan .
Tom hade ingen aning om vad som försiggick .
Tom har en tvillingbror som heter John .
Tom dolde sina bekymmer för sin fru .
Tom leker med sin leksakslastbil .
Tom tycker att Mary är vacker .
Tom vill att Mary ska träffa hans mor .
Tom dömde en konsttävling .
Tom var domare i en konsttävling .
Tom svetsade samman de två rören .
Tom kommer inte att döda någon annan .
Tom undrade varför Mary var så sen .
vi ursäktar avbrottet .
vi måste försöka bryta dödläget .
vi sprang hela vägen till stationen .
vi borde iaktta hastighetsbegränsningen .
vi har en begränsad budget .
vi har varit gifta i fem år .
vad gjorde du i går kväll ?
vad tycker du om att göra på söndagar ?
vad gillar du att göra på söndagar ?
vad tycker du om den här tröjan ?
vad ska du göra på fredag ?
vad ska du göra med den ?
vilken är din favoritprotestsång ?
vilken ordbok syftade du på ?
vilket land är störst , Japan eller England ?
Vilka studerande ska göra provet ?
vilket tåg tänker du ta ?
vem springer snabbast i din klass ?
vem uppfanns telefonen av ?
vem är den där kvinnan i brun jacka ?
varför vill du begå självmord ?
hur kommer det sig att du alltid är sen ?
skulle du vilja ha lite äggröra ?
ni kan välja vilken ni vill .
du borde rensa ogräset .
du blev tillsagd att stanna på skeppet .
du har druckit tre koppar kaffe .
ni har druckit tre koppar kaffe .
&quot; är du svensk ? &quot; &quot; nej , jag är schweizisk &quot; .
en fånge rymde från fängelset .
olyckor av det här slaget sker ofta .
allt du behöver göra är att vänta och se .
Amerika är ett land av invandrare .
tänker du verkligen göra det ?
älskar du mig inte längre ?
först visste jag inte vad jag skulle göra .
först visste jag inte vad jag skulle ta mig till .
kan jag få lite assistans här ?
köpte du den på svarta marknaden ?
förväntade du dig något annat ?
har ni de här skorna i min storlek ?
vet du när Tom kommer tillbaka ?
vet ni när Tom kommer tillbaka ?
behöver du hjälp med att bära något ?
behöver ni hjälp med att bära något ?
förstår du vad du har gjort ?
vill du att jag berättar en historia för dig ?
vill ni att jag berättar en historia för er ?
vill du att jag ska berätta en historia för dig ?
vill ni att jag ska berätta en historia för er ?
vill ni spela tennis med oss ?
Tillåt inte dig själv att bli tjock .
ursäkta mig , jag råkade tappa mina ätpinnar .
Tyskland ligger mitt i Europa .
det tog länge att komma fram till Boston .
Gomorron . dags att vakna .
Godmorgon . det är dags att vakna .
har du läst ut boken ?
har du hittat dina kontaktlinser ?
har du badat än , Takashi ?
han går alltid till jobbet kl. 8.00 .
han frågade mig om jag gillade matematik .
han bad mig kasta tillbaka bollen .
han kopplade på husvagnen på sin bil .
han köpte en ny klänning till sin dotter .
han köpte sin dotter en ny klänning .
han rensade gatan på kastanjer .
han levde inte upp till förväntningarna .
han har dussintals böcker om Japan .
han kliade sig i huvudet av vana .
han skrev ner telefonnumret .
han skrev ned telefonnumret .
han frågar alltid dumma frågor .
han är tre år äldre än hon .
Helsingfors är huvudstad i Finland .
Hallå där ! vad gör du i mitt rum ?
Hallå där ! vad gör ni i mitt rum ?
Hördu ! vad gör du i mitt rum ?
Hörni ! vad gör ni i mitt rum ?
hans hobby är att samla på gamla frimärken .
hur gick det på arbetsintervjun ?
hur mycket tjänar en rörmokare ?
jag är hans vän och kommer så förbli .
jag ser fram emot att träffa dig .
jag är gift och jag har en dotter .
jag är gift och har två barn .
jag väntar på att affärens ska öppna .
jag känner på mig att någonting är fel .
jag står inte ut med det här oljudet längre .
jag kan gå till skolan på tio minuter .
jag går till skolan på tio minuter .
jag kan inte förstå att jag precis sköt mig själv .
jag kan inte fatta att vi äntligen klarade det .
jag kommer inte på hans namn just nu .
jag kunde svära på att någonting rörde sig .
jag förväntar mig inte att du ska vara min vän .
jag vill inte bo i en stor stad .
jag har då aldrig sett på maken .
jag måste lösa problemet på egen hand .
jag vet att pengar inte är allt .
jag lärde mig franska i stället för tyska .
jag må vara galen , men jag är inte dum .
jag spelade tennis med Tom i går .
jag gillar verkligen inte Apple @-@ produkter .
jag säger samma sak om och om igen .
jag borde nog be Tom om ursäkt .
jag känner ännu inte till alla detaljer .
jag studerade en stund i morse .
jag pluggade en stund i morse .
jag trodde Tom vad en fullständig idiot .
jag vill kunna läsa japanska .
jag ville återvända till din by .
jag blev väldigt sårad av dina kommentarer .
jag ska lära dig hur man spelar schack .
jag undrar vart det där skeppet är på väg .
jag undrar vem av er som ljuger .
jag skulle vilja ha en chokladglass .
kan jag få köpa några vykort ?
jag skulle vilja köpa några vykort .
jag skulle inte vilja vara i hennes skor .
jag skulle vilja lägga undan mina ägodelar .
jag är på väg till min systers bröllop .
jag säger bara att möjligheten finns .
jag orkar inte ta mig ned på stan .
jag är ledsen , men jag har ingen växel .
jag har bott sex månader i Kina .
jag har aldrig mått så bra i hela mitt liv .
jag har aldrig sett ett rött kylskåp .
om han ansträngde sig så skulle han lyckas .
Importen av brittiska varor ökade .
det ser ut att bli regn .
alla verkar gilla golf .
det vore trevligt om du kunde komma .
det är ett svårt ord att uttala .
det är en timmes promenad till stationen .
det är inte lätt att lösa problemet .
det är inte viktigt vad jag heter .
Japan är fullt av vackra landskap .
skulle jag kunna få ett glas öl , tack ?
skulle jag kunna få ett glas mjölk , tack ?
skulle jag kunna få ett glas vin , tack ?
det kanske inte kommer att spela någon roll .
det kanske inte spelar någon roll .
män är inte så annorlunda från kvinnor .
min hund låtsas ofta sova .
min pappa går i kyrkan på söndag .
mitt hår är längst i klassen .
min mor sade åt mig att uppföra mig .
min storasyster är bra på att sjunga .
min åsikt skiljer sig från din .
apelsiner innehåller mycket C @-@ vitamin .
vår hund gräver ner ben i trädgården .
vår lärare kommer till skolan med bil .
Papegojor härmar ofta mänskligt tal .
människor agerar inte alltid rationellt .
flytta tv @-@ apparaten till vänster är du snäll .
Säkerheten förhöjdes i staden .
hon kom in helt tårögd .
hon talar inte japanska hemma .
hon pratar inte japanska hemma .
hon har äntligen nått Arktis .
kanske förstår hon senare vad jag menade .
hon klappade sin son på axeln .
hon vill ha en fjärde generationens iPad .
fotboll är populärare än tennis .
det är någonting som gör att dörren inte går upp .
Stockholm är Sveriges huvudstad .
det förklarar varför dörren står öppen .
den ön har tropiskt klimat .
den där röda tröjan ser bra ut på dig .
den där slipsen passar bra till din skjorta .
det är Toms standardsvar .
bebisen sover i vaggan .
pojken gick vilse i skogen .
bron byggdes av romarna .
barnet kastade sten på katten .
matchen blev uppskjuten på grund av regn .
matchen sköts upp på grund av regn .
huset brann ner till grunden .
marken omvandlades till en park .
ju mer vi har desto mer vill vi ha .
flygplanet ankommer klockan åtta .
polisen är här för att tala med dig .
Guldpriset ändras dagligen .
Guldpriset fluktuerar dagligen .
Mötesrapporten är färdig .
tåget avgick i tid .
de två männen var kompanjoner .
det är en massa ägg i lådan .
det finns många parker i London .
det finns inget att klaga på .
det kommer ingenting bra på tv .
det finns yoghurt i kylskåpet .
sådana här saker händer bara i Sverige .
de köpte ett hus på Parkgatan .
de bar in Tom på en bår .
denna byggnad håller på att rasa samman .
det här är en väldigt tidsödande uppgift .
det här är huset som han bor i .
detta är huset han bor i .
det här är vad jag har letat efter .
tre passagerare fick föras till sjukhus .
i dag har jag inte tid för det här .
Tom ser Mary som en hjältinna .
Tom fick inte något gjort idag .
Tom har aldrig ätit rått hästkött .
Tom lär sig att dansa tango .
Tom kan bara inte komma överens med Mary .
Tom skrattade åt alla Marys skämt .
Tom slutade aldrig leta efter Mary .
Tom råkade salta sitt te .
Tom skrattade sällan åt Marys skämt .
Tom fick höra att han var för kort .
Tom var inte som alla de andra pojkarna
Toms mamma gör alla hans kläder .
trafikolyckor sker dagligen .
vi köpte en bit mark tillsammans .
vi kan prata om det i framtiden .
vi har mycket snö vintertid .
vi såg något vitt i mörkret .
vi försökte att kontakta det andra skeppet .
vi kommer att behöva senarelägga mötet .
vi har gäster i morgon kväll .
Vilka djur bebor de där öarna ?
vad ritade han på tavlan ?
vad mer behöver vi prata om ?
vilken är din favoritactionrulle ?
vilken sorts vin rekommenderar du ?
vad är Finlands huvudstad ?
när och var serveras frukost ?
när såg du Tom senast ?
vad föredrar du , Cola eller Pepsi ?
vem var det som faktiskt genomförde operationen ?
varför gjorde du en sådan dum sak ?
varför följer du inte Toms exempel ?
varför följer ni inte Toms exempel ?
varför skulle det spela någon roll ?
Vargar brukar inte attackera människor .
skulle du ha något emot att jag ställer en fråga ?
kan du vara snäll och vänta en minut ?
i går var det söndag , inte lördag .
du och jag har någonting gemensamt .
du kan använda mitt skrivbord om du vill .
det är inte du som bestämmer på det här skeppet .
du måste inte bestämma dig just nu .
det är bäst att du inte väntar längre .
du måste läsa mellan raderna .
man måste läsa mellan raderna .
du passar bra i kort hår .
du måste göra det mycket mer försiktigare .
du måste bli kvitt den där ovanan .
du måste göra dig av med den där ovanan .
du måste sluta ljuga för dig själv .
du borde ha ringt mig med en gång .
du är livrädd , eller hur ?
en katt låg och sov i bastrumman .
en apa klättrar upp för ett högt träd .
en bild säger mer än tusen ord .
alla medborgare borde respektera lagen .
arabiska är ett mycket viktigt språk .
följer du med mig till affären ?
är du alldeles från vettet ?
julen står för dörren .
Columbus upptäckte Amerika 1492 .
kom ner så snart som möjligt .
åt du upp resten av mandlarna ?
satte du på frimärket på brevet ?
har ni några japanska dagstidningar ?
har ni japanska tidningar ?
tror du att vi borde överge skeppet ?
vill du att jag ska hålla ett öga på Tom åt dig ?
vill ni ha te eller kaffe ?
betyder det att du vill göra slut ?
låt inte den här informationen läcka ut .
varje stad i USA har ett bibliotek .
det är fyrtioåtta sjömän på skeppet .
ge henne det här brevet när hon kommer .
han skar ut en buddhastaty ur trä .
han behövde inte ta med sig ett paraply .
han tjänar tre gånger så mycket som jag .
han tjänar tre gånger så mycket som jag gör .
han är alltid villig att hjälpa andra .
han studerade hårt så han inte skulle misslyckas .
han litar mycket på sin assistent .
han anmärkte jämt på mig .
han gick ut en runda med hunden .
han är tillbaks om några dagar .
hennes enda fritidsintresse är att samla på frimärken .
hur hände trafikolyckan ?
hur säger man &quot; adjö &quot; på tyska ?
jag ber om ursäkt om jag har sårat dig .
jag köpte den här kameran för 35 000 yen .
jag kan knappt se utan mina glasögon .
jag kan inte ge dig någonting just nu .
jag kan inte förstå någonting av det han säger .
jag känner inte för att gå ut i kväll .
jag har inget att skriva med .
jag tyckte att den här filmen var väldigt intressant .
jag hade ingen aning om att Tom inte var lycklig här .
jag har en vän som bor i Boston .
jag har en massa arbete att göra imorgon .
jag har ingenting emot förslaget .
jag har inget med brottet att göra .
jag måste åka med min son till läkaren .
jag har inte sett henne sen förra månaden .
jag skrattade väldigt mycket när jag såg det där .
jag lärde mig mycket om grekisk kultur .
jag gillar att gå en tur i parken .
jag gillar den långsamma rytmen i den där sången .
jag tappade bort min väska på väg till skolan .
jag har aldrig problem med att somna .
jag önskar bara att jag kunde hjälpa er alla .
jag beställde boken för över en vecka sedan .
jag utövar yoga utomhus när jag kan .
jag bryr mig verkligen inte om vad Tom tycker .
jag borde ha lyssnat på ditt råd .
jag studerade flitigt när jag gick i skolan .
jag tror Tom letar efter sina nycklar .
jag tror att både Tom och Mary ljuger .
jag trodde att ni två var lika gamla .
det var inte jag som klippte Toms hår .
jag kommer att åka oavsett väder .
jag kommer inte att ha tid med det i morgon .
jag skulle vilja tala med dig igen .
jag skulle vilja tala med er igen .
jag skulle vilja träffa dig igen nästa vecka .
jag vill att du kommer tillbaka nästa vecka .
jag kommer att vara sexton år gammal på min nästa födelsedag .
jag tar ingen semester i år .
jag har aldrig varit hemma hos min farbror .
jag har aldrig varit hemma hos min morbror .
om du inte vill att jag ska åka , så gör jag det inte .
i det här fallet tror jag att han har rätt .
är det okej om jag lånar telefonen ?
finns det något jag kan göra för att hjälpa till ?
det beror på stolens storlek .
det var omöjligt att hitta ett svar .
det var omöjligt att finna ett svar .
det är ingen bra bil , men det är en bil .
Kyoto är känt för sina gamla tempel .
det verkar bli en lång dag i dag .
se till att ingen följer efter dig .
Försäkra dig om att ingen följer efter dig .
kan jag använda telefonen en stund ?
du kanske borde kolla till Tom .
mer än femhundra personer blev skadade .
mer än femhundra personer skadades .
min födelsedag är inte på en månad .
det är en månad till min födelsedag .
det är en månad tills min födelsedag .
min födelsedag är inte förrän om en månad .
min födelsedag är först om en månad .
min bror bor i en liten by .
min pappa tog oss till djurparken i går .
min far varken röker eller dricker .
min pappa jobbar på ett elföretag .
min mormors sjuksköterska är väldigt snäll .
min farmors sjuksköterska är väldigt snäll .
ingen vet säkert hur många människor som dog .
ingen kan göra det så bra som Tom kan .
vår lärare ser ung ut för sin ålder .
lek där ute i stället för att titta på tv .
Religion är ett opium för folket .
hon kan spela den här melodin på piano .
hon ger sin son för mycket pengar .
hon läste hans brev om och om igen .
hon sa att jag borde sluta röka .
hon rörde om i kaffet med en sked .
hon vill hålla honom på avstånd .
hon var tvungen att ge upp planen .
Somliga läser böcker för att slå ihjäl tid .
Vissa läser böcker för att slå ihjäl tid .
Förlåt , jag hade inte med det att göra .
Artikeln var skriven på engelska .
det är väldigt snällt av er att säga det .
Adressen på det här paketet är fel .
stranden var full av turister .
pojken tog tag i kattens svans .
Grannhunden skäller alltid .
bonde plöjde hans fält hela dagen .
Festivalen kommer att gå av stapeln nästa vecka .
det är lätt att ta sig till ön med båt .
den långa resan förvärrade hennes skada .
Romanerna han skrev är intressanta .
Polismannen bär en gasmask .
presidenten har avskaffat slaveriet .
presidenten tillträder sitt ämbete imorgon .
den unga mannen bor i ett gammalt hus .
det är ingen här som heter så .
det var blåsigt den dagen .
de kämpade för religionsfrihet .
de erbjöd gästerna lite kaffe .
de vägrade låta tågen röra på sig .
den här kameran är liten , men mycket bra .
den här ordboken kan komma till användning .
det här är en av Toms favoritböcker .
Tom glömde nästan bort mötet .
Tom kom hit för att be oss om hjälp .
Tom kom hit för att be om vår hjälp .
Tom visste inte var han skulle börja .
Tom diskuterade problemet med Mary .
Tom dricker sex koppar kaffe om dagen .
Tom tar en promenad varje eftermiddag .
Tom har svårt att fatta beslut .
Tom höll upp bildörren åt Mary .
Tom hjälpte Mary att ta av sig jackan .
Tom har dörrarna låsta om natten .
Tom är skyldig Mary trehundra dollar .
Tom satt tyst och tittade på elden .
Tom tycks ha glömt bort mitt namn .
Tom verkar veta vem den där kvinnan är .
Toms tal var rätt underhållande .
Toms tal var rätt så underhållande .
Toms tal var ganska underhållande .
vi kan inte anta att de här pengarna är Toms .
vi kan inte anta att dessa pengar är Toms .
vi kan inte sova på grund av oljudet .
vi hade ett kort lov i februari .
vi gör mjölk till ost och smör .
vi gör ost och smör av mjölk .
vi letar efter en nedgrävd skatt .
vi hinner inte i tid till mötet .
vi ska ha fest på fredag kväll .
vi påverkas av vår omgivning .
vad tycker du att vi ska göra nu ?
det han sa visade sig vara en lögn .
när fick du konsertbiljetten ?
när var första gången du träffade henne ?
vem är flickan som står där borta ?
varför kom du inte hem igår kväll ?
varför kom du inte hem i går kväll ?
väntar du på oss vid stationen ?
väntar du på oss på stationen ?
väntar ni på oss på stationen ?
väntar ni på oss vid stationen ?
kommer du att vänta på oss på stationen ?
kommer du att vänta på oss vid stationen ?
kommer ni att vänta på oss vid stationen ?
kommer ni att vänta på oss på stationen ?
skulle du vilja ha en cappuccino ?
du behöver inte vänta till slutet .
du kan komma med oss om du vill .
du borde ha bett om ursäkt till henne .
du borde köpa en telefonsvarare .
du borde följa skolans regler .
ni borde följa skolans regler .
ni bör följa skolans regler .
du borde tala med din arbetsgivare .
där tar du troligen fel .
det odlas mycket sockerrör på Kuba .
efter måltiden frågade jag efter räkningen .
Al Smiths föräldrar kom från Irland .
Uttalar jag ditt namn korrekt ?
Uttalar jag ert namn korrekt ?
finns det mycket haj här i trakten ?
tänker du ligga i sängen hela dagen , eller ?
tänker du berätta för Tom vad jag gjorde ?
tänker du berätta för Tom vad jag har gjort ?
skynda dig , annars missar du tåget .
skönheten ligger i betraktarens ögon .
morötter och rovor är ätbara rötter .
julen föll på en lördag det året .
det året föll julen på en lördag .
kom igen , jag köper glass åt dig .
skulle jag kunna få ett glas vatten , tack ?
kan du släppa av mig vid biblioteket ?
skulle du kunna upprepa frågan ?
visste du att jag skulle få sparken ?
talade du om för Tom vad Mary hade gjort ?
vet du ens var skolan ligger ?
vet du var mina gamla glasögon är ?
tror du att det kommer att göra någon skillnad ?
tror du det kommer göra någon skillnad ?
tror du att de kan vara farliga ?
gör läxorna innan du tittar på tv .
lägg ingenting på lådan .
det är antingen Tom eller Mary som ljuger .
ta reda på vem Tom har pratat med .
har du redan skrivit på kontraktet ?
har ni redan börjat inreda ?
han frågade mig om jag ville åka utomlands .
han kunde inte komma tillbaka , då han var sjuk .
han tog ett fast tag om tennisracketen .
han hade tre söner som blev advokater .
han har en korg full av jordgubbar .
han är van vid att gå långa sträckor .
han såg ut som om inget hade hänt .
han visade mig hennes fotografi i smyg .
han föddes i en liten stad i Italien .
hennes namn är känt världen över .
hans namn är känt världen över .
hans svar var kort och koncist .
hur kan jag åka buss till sjukhuset ?
hur visste du att jag var kanadensare ?
hur länge tänker du stanna här ?
hur många gånger måste jag säga det till dig ?
jag bad Tom gå och shoppa med Mary .
jag gjorde ett försök att simma över floden .
jag får inte så mycket betalt som jag skulle vilja .
jag vet inte hur man spelar golf överhuvudtaget .
jag vet inte vad det där templet heter .
jag vet inte vad det templet heter .
jag vet inte vad ni vill att jag ska säga .
jag vet inte vad du vill att jag ska säga .
jag vet inte när jag kan ta rast .
jag vet inte varför Tom gjorde som han gjorde .
jag behöver inte höra alla detaljer .
jag förstår inte varför det är en så stor grej .
jag tror inte att det här är Toms paraply .
jag förstår inte vad du håller på med .
jag förväntade mig nästan att Tom skulle börja dansa .
jag har ett tajt schema den här helgen .
jag har inte ätit någonting på sex dagar .
jag har inte ätit på ett par dagar .
jag hoppas att vi har tagit det rätta beslutet .
jag hoppas att vi har tagit rätt beslut .
jag hoppas att vi har fattat rätt beslut .
jag behöver lägga mej ner en stund .
jag behöver bara ligga ner en minut .
jag visste att Tom inte skulle förlora .
jag gillar hundar och min syster gillar katter .
jag tycker om hundar och min syster tycker om katter .
jag älskar naturen , men jag avskyr insekter .
jag gjorde ett allvarligt misstag på provet .
jag begick ett allvarligt misstag på provet .
jag lovade att jag skulle vara tillbaka snart .
jag satte upp en liten koja i trädgården .
jag minns huset som jag växte upp i .
jag pratar med Tom på telefon varje dag .
jag trodde att Tom skulle sova till mitt på dagen .
jag brukar dricka kaffe utan socker .
jag låg på sjukhus i några dagar .
jag låg på sjukhus några dagar .
jag var oförmögen att titta henne i ansiktet .
jag tittade på en svensk film i går kväll .
jag önskar att jag kunde simma lika långt som han .
jag undrar om Tom talar sanning .
jag skulle ha gjort exakt det som du gjorde .
jag skulle ha gjort exakt som du gjorde .
det är fritt för fantasin .
jag är här för att be om ditt samarbete .
på den tiden var jag ännu studerande .
på den tiden gick jag och lade mig tidigare .
det verkar som om du har bestämt dig till slut .
det var Tom som sa att du var sjuk .
det var just likt honom att komma för sent .
det hade inte gjort någon skillnad .
det skulle inte ha gjort någon skillnad .
låt oss sätta upp julgranen här .
Mary är inte Toms biologiska dotter .
min bror har aldrig bestigit Mt Fuji .
min bror är bra på tennis .
min farmor stack iväg med en cowboy .
ingen visste att du var i Tyskland .
en av mina vänner studerar utomlands .
ett , tre och fem är udda tal .
städa golvet med den här moppen , tack .
lägg tillbaka boken där du fann den .
i Europa startar skolorna i september .
hon rådde honom att ta medicinen .
hon förespråkade jämställdhet .
hon blev väldigt arg på barnen .
honom har hon inte sett på länge .
hon har inte sett honom på länge .
hon beordrade honom att städa upp sitt rum .
någon lade ett kuvert på ditt skrivbord .
någon har lagt ett kuvert på ditt skrivbord .
ibland dödas kor av prärievargar .
ibland är det försent att be om ursäkt .
berätta något om ditt land .
allt det hände på bara tre dagar .
orsaken till olyckan är okänd .
kostnaden för boken är fem dollar .
det första steget är det svåraste .
golvet är halt , så var försiktig .
golvet är halt , så var försiktiga .
huset omgavs av en stenmur .
ön träffades av tyfonen .
stegen står i hörnet .
lampan måste fyllas med olja .
polisen har anhållit en misstänkt .
Rosorna blommar i vår trädgård .
affären är öppen året runt .
affären är öppen året om .
ingången till tunnelbanan ligger vid hörnet .
Tunnelbaneingången ligger vid hörnet .
solen sken , men det var ändå kallt .
världen kretsar inte kring dig .
världen kretsar inte kring er .
den här klubben har femtio medlemmar .
du har ett stort hål i strumpan .
det rådde brist på importerad olja .
det fanns nästan ingenting i rummet .
det finns ingen chans att han kommer att återhämta sig .
de här kattungarna är så söta och gosiga .
de lyssnar inte alltid på sina föräldrar .
de lyder inte alltid sina föräldrar .
de gjorde honom till klubbens ordförande .
de säger att han föddes i Tyskland .
det sägs att han föddes i Tyskland .
de bytte plats med varandra .
de kommer att bygga ut sin butik .
den här boken innehåller fyrtio fotografier .
det här är mycket viktigt .
det här är en fråga av stor betydelse .
den här gamla bilen är din om du vill ha den .
denna punkt förtjänar särskild emfas .
det här ägde rum följande dag .
Tom gick med på att åka till Boston med Mary .
Tom höll med om allt som Mary sa .
Tom höll med om allt Mary sa .
Tom bär nästan alltid mörka kläder .
Tom och Mary verkar inte hungriga .
Tom och Mary verkar inte vara hungriga .
Tom och Mary har en tonårig dotter .
Tom och Mary såg lika förvirrade ut .
Tom bad om en filt och en kudde .
Tom frågade om jag skulle vilja laga mat .
Tom frågade mig vad mitt andranamn var .
Tom böjde sig ner och tog upp myntet .
Tom ringde och sa att han skulle bli sen .
Tom kom fram bakom förhänget .
Tom kom fram bakom draperiet .
Tom kan inte tro att Mary är över trettio .
Tom kommer hit så gott som varje dag .
Tom kunde inte höra det , men det kunde Mary .
Tom bestämde sig för att skjuta upp beslutet .
Tom gjorde samma sak som Mary gjorde .
Tom använde inte ordet &quot; omöjligt &quot; .
Tom dog tre veckor efter krocken .
Tom uppskattar inte det som Mary gjorde .
Tom kände sig trött efter att ha jobbat hela dagen .
Tom tvingade Mary att skriva under kontraktet .
Tom tvingade Mary att skriva på kontraktet .
Tom hyste stor kärlek för sitt land .
Tom bjöd in oss till sin sommarstuga .
Tom står inför några allvarliga problem .
Tom är helt enkelt inte så värst bra på att dansa .
Tom är helt enkelt inte särskilt bra på att dansa .
det är Tom som kommer att stå för matlagningen .
Tom är inte min bror . han är min kusin .
Tom ser ut att ha en dålig dag .
Tom måste bestraffas för det som han gjorde .
Tom plöjde sig fram genom folkhopen .
Tom plöjde sig fram genom folkmassan .
Tom tryckte sig fram genom folkhopen .
Tom sätter massor av socker i sitt kaffe .
Tom försvann snabbt in i folkmassan .
Tom sträckte sig efter förstoringsglaset .
Tom sitter bakom Mary på fransklektionerna .
Tom spenderar mycket pengar på kläder .
Tom trodde att Mary kanske inte kände John .
Tom berättade för mig att han var besviken .
Tom sa att de kommer att dö allihop .
Tom sa att alla kommer att dö .
Tom sa att du och Mary dejtade .
Tom gick hastigt genom korridoren .
Tom blev aldrig fälld för brottet .
Tom fälldes aldrig för brottet .
Tom såg sina sondöttrar dansa .
Tom såg sina dotterdöttrar dansa .
Tom kommer aldrig att märka skillnaden .
Toms föräldrar bor i en gammal husvagn .
Toms fru lämnade honom för tre månader sedan .
Vampyrer måste dricka blod för att överleva .
vi såg inga flickor i gruppen .
vi får inte många besökare här nere .
vi hade en fantastisk semester i Sverige .
vi har en reservation klockan halv sju .
vi måste avsluta det här arbetet till varje pris .
vi döpte min son efter min farfar .
vi döpte min son efter min morfar .
vi stötte på dem vid bussterminalen .
vi väntar främmande i kväll .
vi kommer att söka genom hela skeppet .
vi ska söka genom hela skeppet .
vi måste bestämma när vi ska börja .
var det du som ringde polisen ?
vad trodde du att jag skulle göra ?
vad trodde ni att jag skulle göra ?
vad tyckte du om konserten ?
vad exakt är det du tror att Tom gjorde ?
Vilka språk talas i Amerika ?
vilken tid stänger postkontoret ?
vad skulle du göra om du såg ett spöke ?
vad skulle du ha gjort annorlunda ?
vad hade du gjort annorlunda ?
överallt hon kommer är hon uppskattad .
vem röstade du på i valet ?
varför kom du inte hem i går kväll ?
varför avbryter du mig hela tiden ?
kan ni ursäkta mig ett ögonblick bara ?
med Tom hade det varit annorlunda .
går det bra att jag sätter på teven ?
kan ni vänta i några minuter ?
går det bra att ni väntar några minuter ?
i går eftermiddag skrev jag ett brev .
du kan inte klandra henne för vad hon gjorde .
du måste vara en utomordentlig läkare .
du känner antagligen till det som Tom gjorde .
du stötte på honom tidigare , eller hur ?
ni stötte på honom tidigare , eller hur ?
du borde inte ha läst Toms brev .
du borde verkligen inte dricka kranvattnet .
din cykel är mycket nyare än min .
en dag kommer du att få lön för mödan .
&quot; hur gammal är du ? &quot; &quot; jag är sexton år &quot; .
en fladdermus är lika lite fågel som en råtta .
Sedermera antog han en ny identitet .
USA avskaffade slaveriet 1863 .
finns det reserverade platser på tåget ?
Berlin är Tysklands största stad .
kan jag låna ditt suddgummi en stund ?
jämfört med sin far är han ytlig .
såg du verkligen att Tom hjälpte Mary ?
hjälper du alltid Tom att städa sitt rum ?
har du en kofot i verktygslådan ?
kommer du ihåg när du senast såg Tom ?
vill du att jag ber Tom att hjälpa dig ?
gör det ont att ta hål i öronen ?
glöm inte att dricka mycket vatten .
påbörja inte något du inte kan avsluta .
har du skickat in din anmälan än ?
han startar alltid till jobbet kl. 8.00 .
han kände i fickan efter tändaren .
han kände i fickan efter sin tändare .
han gav oss kläder , och pengar också .
han talar jämt illa om sin fru .
han talar alltid illa om sin fru .
han måste köpa en ny cykel åt sin son .
han sa att han skulle åka till Italien .
han sa att han var på väg till Italien .
han besökte ett barnhem i Texas .
han skulle aldrig få se sina föräldrar igen .
han kommer att få veta hemligheten förr eller senare .
han är alltid ivrig att få höra skvaller .
han är vänligt mot alla sina klasskamrater .
hans dumma svar överraskade allihopa .
hans dumma svar överraskade alla .
hur övertygade Tom Mary till att hjälpa oss ?
hur skiljer sig din åsikt från hans ?
hur många äpplen vill du att jag köper ?
hur många äpplen vill du att jag ska köpa ?
hur många äpplen vill ni att jag ska köpa ?
hur många äpplen vill ni att jag köper ?
hur många timmar arbetade du den här veckan ?
hur många människor var ombord på det där skeppet ?
jag kan inte hitta Tom . har han redan gått ?
jag vet ingenting om dinosaurier .
jag vet inte vad som har hänt med honom .
jag tror inte att hon skulle förstå det .
jag vill inte diskutera det med Tom .
jag vill inte veta vad han heter .
jag oroar mig inte så mycket om mitt CV .
jag kände att jag bara var tvungen att komma av skeppet .
jag gav tiggaren alla pengar jag hade .
det hade jag fullständigt glömt bort .
jag åt en halv grapefrukt till frukost .
jag har en vän som klipper sitt eget hår .
jag har en kompis som klipper sitt eget hår .
jag har hört den låten sjungen på franska .
jag har fler kjolar än min storasyster .
jag har inget att göra med det här .
jag måste sätta ett frimärke på kuvertet .
jag hörde att Tom inte sjunger längre .
jag hoppas att din förkylning går över snart .
jag hoppas att du njuter av din vistelse här .
jag hoppas att ni trivs här .
jag vet att jag inte kan kasta boll särskilt bra .
jag vet att jag inte är så duktig på att kasta boll .
jag vet precis vem Tom tänker gifta sig med .
jag tycker om att sjunga och att spela gitarr .
jag tycker om att sjunga och spela gitarr .
jag tycker om att gå och titta på baseboll .
jag föredrar att åka tåg framför att flyga .
jag såg en vit hund hoppa över staketet .
jag skulle ha gått dit själv .
jag borde ha gått dit själv .
jag talar japanska , engelska och franska .
jag pratar japanska , engelska och franska .
jag tycker inte att du borde vänta längre .
jag trodde att Tom skulle säga hej till Mary .
jag ville bli astrofysiker en gång i tiden .
jag ville ringa några telefonsamtal .
jag kommer att förklara detta skämt för dig senare .
jag ska ta med dig till mitt palats imorgon .
jag ska ta med er till mitt palats imorgon .
jag är trött på att äta på restaurang .
jag lyssnar på Björks senaste låt .
jag är inte det minsta intresserad av kemi .
jag har känt Tom sedan vi var barn .
jag har känt Tom sen vi var barn .
om man äter för mycket blir man tjock .
om du äter för mycket kommer du att bli tjock .
vilket år föll Berlinmuren ?
är Tom fortfarande kapten över ditt skepp ?
det måste inte göras nu med en gång .
det låter som om du faktiskt menar det .
man trodde att valar var fiskar .
titta på den där byggnaden . är det ett tempel ?
vi borde kanske prata om det här först .
mamma var allt som oftast väldigt upptagen .
min bror har aldrig bestigit Mt Fuji .
min bror måste skriva en tentamen .
mitt huvudämne är europeisk medeltidshistoria .
min mor tar en tupplur varje eftermiddag .
mina föräldrar dog när jag var mycket ung .
min föraning visade sig vara rätt .
en gång i tiden trodde man att människor inte kunde flyga .
Osmanska turkar erövrade Egypten år 1517 .
vårt skepp blev inte skadat i striden .
hon hjälpte den gamla mannen över vägen .
hon läser tidningen varje morgon .
hon ville gifta sig omedelbart .
hon bar babyn på ryggen .
tala högre så att alla kan höra dig .
tennis är väldigt populärt bland studerande .
det är ett av mina favorituttryck .
flygplanet lyfte för tio minuter sedan .
Fåglarna flög iväg åt alla håll .
företaget vill anställa 20 personer .
hissen verkar vara trasig .
fienden förstörde många av våra skepp .
ön är ett paradis för barn .
Juvelen stals under natten .
polisen arresterade honom för smuggling .
Prinsessan låg och blundade .
Trottoarerna var blöta efter regnet .
New Yorks gator är väldigt breda .
läraren välkomnade de nya studenterna .
Tornet lutade lätt till vänster .
staden förstördes under kriget .
det finns nästan inget syre i rummet .
det fanns några barn i rummet .
det var några barn i rummet .
det är ingen på det här skeppet förutom oss .
det finns inte plats för alla .
de är nöjda med det nya huset .
de är väldigt intresserade av astronomi .
de hämtar våra sopor varje måndag .
de förklarade sig oskyldiga .
de var medlemmar av medelklassen .
det här är mannen som jag letat efter .
den här gamla bilen går sönder hela tiden .
Tom valde att inte kommentera saken .
Tom ville inte gå dit med Mary .
Tom ville inte åka dit med Mary .
Tom tycker inte om huset han bor i .
Tom vet inte om att jag är Marys pojkvän .
Tom vet inte att jag är Marys pojkvän .
Tom tycker inte om att prata om sport .
Tom gillar inte att prata om sport .
Tom är förväntad att anlända inom kort .
Tom är ute på gården och räfsar löv .
Tom är van att ta snabba beslut .
Tom är inte den gitarrist som han brukade vara .
Tom ser ganska mycket äldre ut än Mary .
Tom rörde sig genom den svagt upplysta gränden .
Tom insåg att Mary hade något i kikaren .
Tom insåg att Mary hade något fuffens för sig .
Tom insåg att Mary hade något för sig .
Tom säger att han inte har någon aning om var Mary är .
Tom säger att han inte har en aning om var Mary är .
Tom sade till Mary att hålla dörren stängd .
Tom sade åt Mary att hålla dörren stängd .
Tom önskar att han inte hade gjort det han gjorde .
Tom kommer inte , och inte Mary heller .
Tom skulle aldrig döda sin egen dotter .
Toms mamma glömde att packa ner hans lunch .
Toms party var ganska roligt , faktiskt .
Toms självmord ändrar ingenting .
två barn sitter på staketet .
två personer kommer in på den här biljetten .
vi behöver faktiskt inte göra det nu .
så här kan vi inte fortsätta länge till .
vad ska du göra ikväll ?
vad hände med resten av maten ?
hur mycket förbrukar den här bilen ?
hur dags gick du och lade dig i går ?
var är fjärrkontrollen till tv:n ?
skulle du vilja äta lunch tillsammans ?
skulle du kunna sänka radion ?
du gjorde rätt som berättade för oss .
du måste inte komma hit varje dag .
du ser precis ut som din storebror .
du påminner om en pojke som jag kände .
du ville att det skulle bli så här , eller hur ?
många människor dödades i kriget .
en ung flicka satt vid ratten .
alla dörrar i huset var stängda .
allt du behöver göra är att trycka på knappen .
vilken blomma som helst går bra , så länge den är röd .
finns det några biografer här i närheten ?
pojkar härmar ofta sina idrottshjältar .
men det var förstås länge sedan .
skulle jag kunna få prata med dig en stund ?
kan du sänka priset till tio dollar ?
kan du skriva ut det här dokumentet åt mig ?
barn behöver en lycklig hemmiljö .
lektionen börjar inte förrän halv nio .
kom tidigt så vi kan diskutera planerna .
skulle ni barn kunna hjälpa mig att duka av bordet ?
Demokratin har sitt ursprung i antikens Grekland .
Detroit är känt för sin bilindustri .
sa Tom hur länge han skulle vara i Boston ?
hittade du det du sökte efter ?
gillar du glass med kinuskismak ?
tror du att vi kommer att hitta hennes hus ?
tror ni att vi kommer att hitta hennes hus ?
tror du att du kommer att kunna hjälpa mig ?
kommer Tom bra överens med andra människor ?
förstår du dig på den här rapporten ?
glöm inte festen nästa vecka .
glöm inte att det finns undantag .
vet du inte vad som hände i går ?
har du skrivit upp telefonnumret ?
har du skrivit ned telefonnumret ?
han kan inte ha sagt något så dumt .
han inser inte att han är tondöv .
han förklarade varför experimentet misslyckades .
han bröt nacken i olyckan .
han gick vilse när han var ute och gick i skogen .
han har alltid hängivit sig åt musik .
han har god anledning att tro det .
han anmärker jämt på andra .
han lider av en svår sjukdom .
han kysste sin dotter på pannan .
han gick ut ur rummet utan att säga ett ord .
där såg han det han hade drömt om .
han visade mig en massa vackra bilder .
han visade mig massor av vackra bilder .
han vill spela fotboll i eftermiddag .
han gick ut trots ösregnet .
han klagar alltid på maten .
hans bok blev föremål för kritik .
hans otrevliga kommentarer spädde på dispyten .
hur tidigt går du upp om morgnarna ?
hur långt borta tror du att det där skeppet är ?
hur många språk finns det i Europa ?
hur många moskéer finns det i Istanbul ?
jag är finsk , men jag talar svenska också .
jag kommer att gå av vid nästa hållplats .
jag ville inte säga det till dig på telefon .
jag har inga rena kläder att använda .
jag vet inte exakt när jag kommer att komma tillbaka .
jag vet inte vad han är för slags person .
jag vet inte var jag har lagt min mobiltelefon .
jag vet inte varför Tom behövde göra det .
jag schamponerar inte håret på morgonen .
jag tvättar inte håret på morgonen .
jag tror inte att Tom gjorde någonting med den .
jag tror inte att Tom gjorde någonting med det .
jag tror inte att Tom gjorde något med det .
jag tror inte att Tom talar sanning .
jag tror inte Tom vet hur man gör det .
jag tror inte att Tom var berusad .
det tycker jag inte är en särskilt bra idé .
jag tycker om att titta på gamla familjebilder .
jag lärde känna honom när jag var student .
jag har inte pratat med Tom om det än .
jag hoppas att jag inte behöver använda den här pistolen .
jag hoppas att vi ses igen snart .
jag hoppas att vi ses snart igen .
jag måste få det färdigt så fort som möjligt .
jag spelade ofta fotboll när jag var ung .
jag måste ändå fråga Tom om lov .
jag tror att Tom inte förstod skämtet .
jag trodde aldrig att Tom skulle sluta prata .
jag översatte dikten så gott som jag kunde .
jag vill spela tennis med dig någon dag .
jag vill spela tennis med dig någon gång .
jag vill att du överger den här dumma planen .
jag var i Boston med frugan i förra veckan .
jag ska fråga honom om det imorgon då .
jag skulle vilja boka ett flyg till Vancouver .
jag skulle vilja följa med , men jag är pank .
jag är riktigt oroad över din framtid .
du kommer säkert på nånting .
det spelar ingen roll längre .
det hände att hon tog ett bad .
det är omöjligt att leva utan vatten .
det är inte döden jag fruktar , utan att dö .
det ser ut som att alla från byn är här .
det tog en månad för min förkylning att gå över .
det var en väldigt svår historia att skriva .
det var hans tystnad som gjorde henne arg .
det skulle inte spela någon roll ändå .
det är viktigt att du berättar sanningen .
det är viktigt att följa en sträng diet .
January är årets första månad .
förra veckan var jag i Boston med min fru .
många använder uttagsautomater för att ta ut pengar .
de flesta japanska tempel är gjorda av trä .
min far är på promenad i parken .
min fru och jag kom överens om en semesterplan .
att spela tennis är bra för hälsan .
snälla fråga inte en sådan fråga .
hjälp mig att översätta det här dokumentet , tack .
kaniner har långa öron och korta svansar .
tomten stod på tomten .
hon slog ihjäl honom med en golfklubba .
hon kunde inte komma för hon var sjuk .
hon försökte inte att översätta brevet .
hon antydde att hon kanske skulle studera utomlands .
hon är en svår person att ha och göra med .
hon lever på grönsaker och råris .
hon stod upp och gick mot fönstret .
hon vill veta vem det var som skickade blommorna .
hon går ofta och shoppar på helger .
Solenergi är en ny energikälla .
en del fabriker förorenar miljön .
förr eller senare kommer sanningen fram .
sluta klaga och gör som du blivit tillsagd .
säg till alla att jag är allergisk mot jordnötter .
Golden Gate @-@ bron är gjord av järn .
Äppelträdet har en vacker blomning .
pojken tömde tallriken på ett ögonblick .
byggnaden uppe på kullen är vår skola .
byggnaden som jag såg var väldigt stor .
Brevets innehåll var hemligt .
dagarna blir allt längre .
läkaren kom i grevens tid .
hunden har bitit hål på min ärm .
dörrarna var låsta utifrån .
Misslyckandet beror på hans vårdslöshet .
gisslan släpps fri imorgon .
gisslan kommer att släppas i morgon .
Advokaten förklarade den nya lagen för oss .
vädret har varit dåligt i två veckor .
deras varor är av högsta kvalitet .
det finns många typsnitt att välja bland .
det var många människor i rummet .
de är som dag och natt .
de efterlyste ett slut på striderna .
de bor i ett nytt hus nära parken .
det här är en bild på skeppet som jag var på .
det här är huset , i vilket min farbror bor .
det här är huset som min farbror bor i .
den här romanen är översatt från engelska .
det här stället har en mystisk atmosfär .
till min förvåning var han bra på att sjunga .
Tom kom faktiskt på det själv .
Tom och Mary fick ändra planerna .
Tom trodde på allt som Maria sa .
Tom kunde inte tro på det som hänt .
Tom ville inte gå dit efter mörkrets inbrott .
Tom ville inte åka dit efter mörkrets inbrott .
Tom delade tårtan i åtta bitar .
Tom pratar faktiskt inte mycket Franska .
Tom kan inte spela piano .
Tom arbetar inte lika hårt som han brukade .
Tom är en ganska bra korgbollsspelare .
Tom kör aldrig för fort .
Tom håller alltid hastighetsbegränsningen .
Tom tog fram sitt häfte och sin penna .
Tom tog fram sitt häfte och sin blyertspenna .
Tom sköljde schampot ur håret .
Tom sade att han tyckte att jag verkade imponerad .
Tom borde ha följt Marys råd .
Tom visade Mary hur man gör det rätt .
Tom tog av örngottet från kudden .
Tom vill att hans pappa köper en ponny till honom .
Toms cykel blev stulen av en narkoman .
Toms cykel blev stulen av en knarkare .
Toms gammelmorfar föddes blind .
Toms gammelfarfar föddes blind .
vi frågar läraren frågor varje dag .
vi hinner med tåget .
vi gillade maten , speciellt fisken .
vi gick ut på en promenad efter frukost .
vi har haft fint väder en tid nu .
vad krävs för att man ska få lite hjälp ?
vad har du där i din ficka ?
vilken sorts spel tycker du om att spela ?
vilken tunnelbanelinje går till stadskärnan ?
vilken tunnelbanelinje går till centrum ?
vilken Harry Potter @-@ bok är din favorit ?
när lämnar din far sitt kontor ?
var var du när jag behövde din hjälp ?
vem har sagt att Tom och jag dejtar ?
varför finns det ingen fisk i den här dammen ?
du är en ängel som handlar åt mig .
du står näst på tur för en befordran .
du kan använda ett lexikon till den här tentamen .
du kan välja vilken bok du vill .
ni får välja vilken bok som helst .
du måste sätta mer vatten i vasen .
du frågar ofta frågor som jag inte kan svara på .
du lovade mig att du skulle ta hand om Tom .
du låg och sov när jag kom hem .
du har förlorat koncentrationsförmågan .
plötsligt blev det mulet .
kommer du någonsin gifta dig igen ?
men vad gör du om han inte kommer ?
kan någon förklara detta för mej ?
äter du kött eller är du vegetarian ?
äter ni kött eller är ni vegetarianer ?
har du en gräsklippare jag kunde låna ?
vill du att jag ska berätta vad Tom gjorde ?
vill du att jag ska berätta för dig vad Tom gjorde ?
är det någon som vet var jag kunde hitta en sådan ?
vet någon var jag kunde hitta en sådan ?
glöm inte att vi måste göra läxorna .
allting var förberett långt i förväg .
har du kollat oljenivån nyligen ?
har du någonsin haft de här symtomen tidigare ?
han kände sig obekväm i sin fars närvaro .
han har vattnet rinnandes i badkaret .
han håller jämt på och styr och ställer .
han verkade besviken över resultaten .
han skrev en bok om djungeläventyr .
han är väldigt smart , så alla gillar honom .
hennes storasyster gifte sig förra månaden .
hur länge ska du vara i Japan ?
jag är hungrig för jag har inte ätit lunch .
jag kan inte fatta att Tom kan teckenspråk .
jag kan inte läsa franska , och ännu mindre tala det .
jag kan inte läsa franska , inte heller kan jag tala det .
jag kan inte säga exakt var problemet är .
jag känner inte för att äta någonting idag .
jag vet inte vad rätt svar är .
jag läser inte lika mycket böcker som jag gjorde tidigare .
jag vill inte prata om det just nu .
jag köpte en ny hatt på köpcentret .
jag hade en bra anledning att inte vara där .
jag har en känsla av att hon kommer att komma idag .
jag har ingen aning om vad Tom pratar om .
jag har spenderat mycket pengar på mitt hus .
jag hörde just vad som hände med Tom .
jag vet precis vad Tom kommer att säga .
jag fick dig att känna dig obekväm , inte sant ?
jag måste göra klart läxan innan middagen .
jag förstod aldrig riktigt vad som hände .
jag sade aldrig att det inte var en bra idé .
jag sa aldrig att det inte var en bra idé .
jag lade märke till att hon satt på första raden .
jag svär att jag aldrig ska göra det igen .
jag tror att vi har köpt allt som vi behöver .
jag tycker att din engelska har blivit mycket bättre .
jag tror inte att din teori håller .
jag tänkte att jag kanske kan köpa dig en drink .
jag trodde att du hade en överenskommelse med Tom .
jag vill ha två korv med bröd med mycket peppar .
jag var irriterad över att hon fortfarande sov .
jag gick och lade mig lite senare än vanligt .
jag lämnar tillbaka boken så fort jag kan .
jag skrev till honom av en helt annan anledning .
jag skulle vilja ha ert svar med en gång .
jag ser fram emot sommarlovet .
Förlåt , det var inte min mening att sparka dig .
jag är ledsen , men det finns ingenting jag kan göra .
jag har alltid varit intresserad av politik .
finns det en tvättmaskin i huset ?
det är länge sedan jag såg honom .
det är en sjukdom som inte kan förebyggas .
det verkar som att du inte tar mig på allvar .
det verkar som att ni inte tar mig på allvar .
det tog mig tre dagar att läsa den här boken .
man trodde att jorden var platt .
det var lättare att göra än jag hade tänkt mig .
det är svårt att förstå hans teori .
nästan allt som Tom säger är lögn .
många vackra blommor blommar på våren .
många turister kommer för att se vattenfallet .
miljoner vilda djur lever i Alaska .
min farfar hör lite dåligt .
min morfar hör lite dåligt .
mitt skosnöre fastnade i rulltrappan .
vår bil är tre år äldre än er .
vår bil är tre år äldre än din .
vår bil är tre år äldre än era .
vår bil är tre år äldre än dina .
snälla rätta mig när jag gör fel .
snälla gå ut ur mitt kontor genast .
Hajfenssoppa är väldigt populärt i Kina .
hon blev tvungen att förlita sig på sin inre styrka .
hon vet bättre än att argumentera med honom .
hon hjälpte dem med bagaget .
hon älskar att se på tennismatcher på tv .
hon älskar att titta på tennismatcher på tv .
hon borde ha gjort klart sina läxor .
hon räckte upp handen för att få bussen att stanna .
hon kommer att bli glad när hon förlovar sig .
Konstiga saker hände på hennes födelsedag .
Konstiga saker skedde på hennes födelsedag .
tv hjälper oss att bredda vår kunskap .
det har gått tio år sedan jag kom hit .
Texas är nästan dubbelt så stort som Japan .
det besegrade laget lämnade så sakta planen .
Diamanten värderades till 5 000 dollar .
Juryn fann mannen skyldig till mord .
månen är mycket vacker i kväll .
soldaterna var utrustade med vapen .
problemet med honom är att han är lat .
det finns knappast några böcker i detta rum .
det finns många galaxer i universum .
det finns bara tre tjejer i klassen .
det ligger en sax på bordet .
det låg nånting på marken .
de blev fördröjda på grund av kraftigt snöfall .
den här boken finns bara tillgänglig i en affär .
det här är Carrie Underwoods senaste album .
det här är det bästa skepp som jag någonsin varit på .
den här kniven är för slö för att skära med .
Tom fick faktiskt Mary till att dansa med honom .
Tom håller med om mycket av det som Mary sa .
Tom dricker alltid kaffe på morgonen .
Tom tror att Mary fattade rätt beslut .
Tom kan tala tre olika språk .
Tom känner inte att han kan lita på Mary .
Tom tror inte att detta är någon tillfällighet .
Tom är förlovad med Marys lillasyster .
Tom sjunger ofta när han är i duschen .
Tom pratar bara franska med sina föräldrar .
Tom sa att han läste en bok om det här skeppet .
Tom pratar bara franska med sina föräldrar .
Tom satt mer än tre år i fängelse .
Tom spenderade mer än tre år i fängelse .
Tom satt mer än tre år i fängelset .
Tom satt över tre år i fängelset .
Tom sov över hos en kompis .
Tom brukade hata Mary . nu älskar han henne .
Tom talar om det för dig när han känner för det .
Tom undrade om det som Mary sade var sant .
vi insåg inte att vi var så högljudda .
natten är ju ganska lång , eller hur ?
hur dags gick du och lade dig igår ?
hur dags gick du och lade dig i går ?
vilket är ditt favoritprogram på tv ?
när katten är borta dansar råttorna på bordet .
vilken tycker du bäst om , Cola eller Pepsi ?
varför måste alla lära sig engelska ?
stör det dig om jag sätter på tv:n ?
skulle du vilja spela tennis på söndag ?
skulle du inte vilja ta lite frisk luft ?
skulle du inte hellre göra det själv ?
du behöver inte gömma någonting för mej .
du klagar så gott som aldrig på någonting .
ni klagar så gott som aldrig på någonting .
för länge sedan fanns det en bro här .
det bodde en vild folkstam där på den tiden .
en liten vinst är bättre än en stor förlust .
det är fritt inträde under jullovet .
alla Toms kläder är gjorda av hans mamma .
Pojkband var mycket populära vid den tiden .
Pojkband var mycket populära på den tiden .
kan du säga namnet på alla träd i trädgården ?
visste du inte att det här skulle hända ?
lova mig att du inte gör det .
han blåste på sina fingrar för att värma dem .
han stannade upp mitt sitt anförande .
han har inga vänner att leka med .
han gick in på banken utklädd som en vakt .
han fick sitt vänstra ben skadat i en olycka .
han är en av Spaniens mest kända författare .
han gick ut ur rummet så fort som jag gick in .
han övertalade sin fru att inte skilja sig .
han skrev ner sina tankar i sin anteckningsbok .
han verkade trivas med sitt liv och sitt arbete .
han stoppade näsduken i fickan .
han mötte några svårigheter .
han gick till affären för att köpa lite apelsiner .
han kommer inte att stanna mer är fyra dagar .
han kommer inte att stanna i mer än fyra dagar .
hej . det är du som är Tom va ? det var längesen .
hans far vigde sitt liv åt vetenskapen .
hans översättning ligger nära originalet .
hur lärde du dig att spela fiol ?
hur länge kommer det här kalla vädret att fortsätta ?
hur ofta byter du rakblad ?
jag har alltid en ordbok nära till hands .
jag antar att du är beredd att ta risken .
jag tror att han kommer att bli rik en dag .
jag står inte ut med oljudet längre .
jag kan inte komma ihåg den låtens melodi .
jag trodde inte att Tom faktiskt skulle prova det .
jag vet inte exakt när jag kommer att vara tillbaka .
jag tycker inte om när du tar med dig jobb hem .
jag gillar inte kvinnor utan personalitet .
jag tror inte att det kommer att regna i morgon .
jag tror inte det finns en doktor här
det känns som om jag sett den här filmen förut .
det känns som om jag har sett den här filmen förut .
jag har ingen aning om vad Tom pratar om .
jag vet att du inte ville att Tom skulle åka in i fängelse .
mitt huvudämne på universitetet var kemi .
jag missade tåget med bara några minuter .
jag tror att Tom och John är enäggstvillingar .
jag tycker att det är tragiskt att inte ha några vänner .
jag tycker att du borde komma och stanna hos mig .
jag trodde att Tom skulle stanna lite längre .
jag vill äta något som inte är sött .
jag vill äta någonting som inte är sött .
jag var väldigt trött , så jag gick och la mig tidigt .
jag var väldigt trött , så jag gick och lade mig tidigt .
jag skulle vilja ställa dig några till frågor .
jag skulle vilja att du betalar i förskott .
jag ska bara ta en promenad för att rensa huvudet .
jag är ledsen , jag tror inte att jag kommer kunna .
jag är förvånad att han antog erbjudandet .
jag är förvånad att han accepterade erbjudandet .
jag är mycket glad att lära känna er .
jag har sett fram emot att få träffa dig .
hade jag vetat skulle jag ha sagt det till dig .
om du vill ta en paus , så säg bara till .
vi råkade befinna oss på samma buss .
det vore bra om vi kunde träffas igen .
det vore kul om vi kunde träffas igen .
hon är kvart över nio .
av ren nyfikenhet , vad skulle du göra ?
många ryssar krävde ett slut på kriget .
kan jag få ett par ostsmörgåsar ?
skulle jag kunna få ett par ostsmörgåsar ?
ingen vet om han älskar henne eller inte .
ingen vet vare sig han älskar henne eller inte .
inte en människa syntes till i byn .
spring fort , annars kommer du för sent till skolan !
ibland vill man bara äta choklad .
sådant kan hända då och då .
det var i det huset som jag föddes i .
olyckan berodde på vårdslös körning .
företaget gör reklam för en ny bil på tv .
företaget marknadsför en ny bil på tv .
Föraren vred ratten åt höger .
Gorillan var ett år gammal vid det tillfället .
huset höll på att målas av min far .
ju mer pengar vi har , desto mer vill vi ha .
nästa konsert kommer att hållas i juni .
den nuvarande regeringen har många problem .
det värsta med sommaren är värmen .
det fanns en lista på tillgängliga kandidater .
det var en massa möbler i rummet .
det var femtio passagerare på planet .
det finns nästan ingen mjölk kvar i glaset .
ett bra vin behöver inte annonseras .
de bor i en liten by i England .
den här klänningen kan se lustig ut , men jag gillar den .
det här är ett postkontor och det där är en bank .
den här stenen är dubbelt så tung som den där .
det här ordet betyder flera olika saker .
till min förvåning så hade han en vacker röst .
Tom visade upp innehållet i sin plånbok .
Tom kommer inte överens med sina grannar .
Tom samlade ihop alla sina saker .
Tom var tolv när Berlinmuren föll .
Tom undrade vad Mary skulle säga till John .
vi klarar oss utan tv , eller hur ?
vi kan se tusentals stjärnor på himlen .
vi vill inte skrämma bort barnen .
vi hade många bra stunder i vår husbil .
när jag öppnade dörren hade jag sönder låset .
när var senaste gången Tom pratade med dig ?
vart går du oftast och klipper dig ?
vem vikarierar för Tom medan han är borta ?
varför är du inte redan ombord på skeppet ?
varför plockar du aldrig undan efter dig ?
skulle du kunna förklara reglerna för mig , tack ?
skulle ni kunna förklara reglerna för mig , tack ?
man behöver kramsnö för att göra bra snöbollar .
man bör alltid tänka innan man talar .
du borde vara försiktigare nästa gång .
du borde vara noggrannare nästa gång .
ni borde vara noggrannare nästa gång .
du måste ta tjuren vid hornen !
din attityd gentemot kvinnor är stötande .
ditt namn har tagits bort från listan .
under förra året skedde det många trafikolyckor .
många tror att fladdermöss är fåglar ..
många människor tror att fladdermöss är fåglar .
en man kom fram till mig och bad om en tändsticka .
Luftföroreningar är ett allvarligt globalt problem .
tror du på spöken ?
känner du mannen som pratade med mig ?
minns du den gången vi åkte till Paris ?
oroa dig inte . han förstår inte tyska .
varje familj har ett skelett i garderoben .
alla vill träffa dig . du är känd !
allt måste handskas med väldigt försiktigt .
var snäll och ge oss två knivar och fyra gafflar .
Hawaii har fint väder året runt .
han gör ingenting annat än klagar dagarna i ända .
han tog sitt liv genom att hoppa ner från en bro .
han tjänar tre gånger så mycket pengar som jag gör .
han tjänar tre gånger så mycket pengar som jag .
han anklagades för att ha stulit dinosaurieben .
hans frånvaro igår berodde på förkylning .
hur många syskon har du ?
jag minns inte exakt vem som sa det till mig .
jag minns inte exakt vem som sade det till mig .
jag kommer inte ihåg exakt vem som sa det till mig .
jag kommer inte ihåg exakt vem som sade det till mig .
jag glömde att klistra på ett frimärke på kuvertet .
jag har inte skrivit ett brev på länge .
jag vet att du gör så bara för att reta mig .
jag gav tillbaka kniven som jag hade lånat .
jag såg dem alla åtta för ungefär en timme sedan .
jag tror att det är dags för mig att skaffa ett nytt jobb .
jag tror att vi har köpt allt som vi behöver .
jag tycker att du borde tänka på framtiden .
jag tycker att du är lite för försiktig .
jag tror att du är lite för försiktig .
jag tycker att du är lite för noggrann .
jag tror att du är lite för noggrann .
jag tyckte jag sa åt dig att inte stå i vägen för mig .
jag trodde att polisen letade efter Tom .
jag var nära att dö av en hjärtattack .
jag höll på att titta på tv när telefonen ringde .
jag tittade på tv när telefonen ringde .
jag kunde inte gå på hans födelsedagskalas .
jag åkte på en tiodagarsresa till Påskön .
jag önskar att jag inte behövde jobba den här helgen .
jag undrar varför hon inte berättade om det för honom .
jag ska plugga engelska i eftermiddag .
jag ska studera engelska i eftermiddag .
jag är van vid att dricka kaffe utan socker .
om jag vore du , skulle jag lyssna på Toms råd .
är det faktiskt så ohälsosamt att äta äggulor ?
det är inte lönt att försöka lösa det här problemet .
det är ingen mening med att försöka lösa det här problemet .
det är inte säkert att köra bil utan bilbälte .
det tog dem två år att bygga huset .
det var svårt för dem att ta sig till ön .
det dröjer inte länge innan hon är tillbaka .
det är kallt , så jag vill äta någonting varmt .
det är knappast värt att bry sig om honom .
det är varmt , så jag vill äta någonting kallt .
det är första min far skrev .
det är dags för dig att sluta titta på tv .
se till att Tom håller sig borta från min dotter .
Mary var Toms flickvän för ett par år sedan .
mor stannade i bilen medan far handlade .
mamma stannade i bilen medan pappa handlade .
de flesta slott omges av en vallgrav .
mor köpte två flaskor apelsinjuice .
min väckarklocka ringde inte i morse .
min far har slutat röka på grund av sin hälsa .
ingen av eleverna var sen till skolan .
snälla , lova mig att du inte gör om det där .
hon frågade var huset låg .
hon vann första pris i en matätartävling .
hon gifte sig mot sin fars vilja .
hon har en ödletatuering på låret .
hon är väldigt duktig på att imitera sin lärare .
hon lyckades avsluta arbetet själv .
hon valde en hatt som matchade hennes klänning .
hon är för ung för att skaffa körkort .
Vissa fiskar kan byta kön .
Publiken bestod mest av elever .
barnet tigger alltid om någonting .
Följden blev att hon förlorade jobbet .
Bristen på pengar är roten till allt ont .
det enda språk Tom kan tala är franska .
det enda språk som Tom kan tala är franska .
polisen lyckades hitta brottslingen .
stadens snabba tillväxt överraskade oss .
vädret är sämre i dag än i går .
hela familjen hjälpte till med att skörda vetet .
det finns en park i centrum .
det är någonting med honom som jag inte tycker om .
det låg glasskärvor över hela golvet .
det fanns inga tecken på liv på ön .
det finns två hundra personer i rummet .
det kommer att finnas mycket tid till det senare .
det kommer det att finnas mycket tid till senare .
det kommer att finnas mycket tid för det senare .
det kommer det att finnas mycket tid för senare .
de skyndade sig till olycksplatsen .
de såg antagligen vårt skepp komma in i hamnen .
de stödde honom och hans politik fortfarande .
det här är bilden som jag tog på Toms hus .
det här är templet som vi brukade besöka .
Tofu kan användas som ersättning för kött .
Tom gjorde faktiskt det han sa att han skulle göra .
Tom gick med på att hjälpa Mary städa köket .
Tom klagar nästan aldrig på någonting .
Tom behöver sannerligen inte mer pengar .
Tom förstår inte vad du säger .
Tom använder tandtråd minst en gång om dagen .
Tom har aldrig klippt sina egna barns hår .
Tom kan komma på vår fest i morgon .
Tom tycker om att lyssna på gamla radioprogram .
Tom gör världens bästa spagetti .
Tom gör världens bästa spaghetti .
Tom masserar tinningarna med sina fingrar .
Tom visade mig brevet som han fick av Mary .
vi kan inte vara utan vatten ens för en dag .
vi kunde inte gå ut på grund av tyfonen .
vi glömde att ta det i beaktande .
vi hade roligt på stranden igår .
vi hade roligt på stranden i går .
vi måste försvara vårt land till varje pris .
vi känner till fler än 100 miljarder galaxer .
vi ska presentera idén för kommittén .
vi ska presentera idén för utskottet .
vi ska se en utländsk film ikväll .
var du nervös under arbetsintervjun ?
vad fattas dig ? du ser blek ut .
vilken är din favoritsnabbmatsrestaurang ?
varför frågar du inte din lärare om råd ?
man kan lära sig många ord genom att läsa .
man kan inte stoppa tillbaka tandkräm i tuben .
du ser ut som en liten flicka i den klänningen .
man stöter på japanska turister överallt .
&quot; skicka mig saltet , tack &quot; . &quot; Varsågod &quot; .
&quot; vad är det där ? &quot; &quot; hur ska jag veta ? &quot;
&quot; vad är det där ? &quot; &quot; hur ska jag kunna veta ? &quot;
en japansk trädgård har vanligtvis en damm .
ett ögonblicks tvekan kan kosta en pilot livet .
var alltid smartare än de personer som anställer dig .
kan du tro att detta faktiskt händer ?
kan du kolla om telefonen är trasig ?
Barnaga är förbjudet i Sverige .
var det svårt att hitta ?
skrev du något i din dagbok idag ?
varje del av ön har utforskats .
att bli klar med detta jobbet innan tisdag kommer att vara enkelt .
att blir klar med det här jobbet innan tisdag kommer att bli enkelt .
att bli klar med det här jobbet innan tisdag kommer att vara enkelt .
att bli klar med detta jobb innan tisdag kommer att bli enkelt .
att bli klar med detta jobb innan tisdag kommer att vara enkelt .
har du skrivit klart din uppsats ?
han stoltserar alltid med sina engelskkunskaper .
han får göra vad han vill med pengarna .
han kan göra vad han vill med pengarna .
han utförde arbetet så gott han förmådde .
han har en chans att tangera det gamla rekordet .
han har inte bytt kläder på två veckor .
han vande sig kvickt vid det kalla vädret .
han vande sig snart vid det kalla vädret .
han använde hennes cykel utan att fråga om lov .
han gick långsamt så att barnet kunde följa med .
han gick långsamt så att barnet kunde hänga med .
han gick långsamt så att barnet kunde hinna med .
han gick sakta så att barnet kunde hinna med .
han gick sakta så att barnet kunde hänga med .
han gick sakta så att barnet kunde följa med .
hur mycket kostar två honungsmunkar ?
jag kan inte tacka nog för din vänlighet .
jag tror inte att det kommer att regna i eftermiddag .
jag tycker inte att den här fåtöljen är bekväm .
jag kände mig väldigt lättad när jag hörde nyheten .
jag hoppas att du kommer fram med en bättre plan .
jag vet att Mary är vackrare än jag .
jag vet att Mary är vackrare än mig .
jag behöver en blyertspenna . kan jag låna en av dina pennor ?
jag vill verkligen veta vad det är som pågår här .
jag har fortfarande inte funnit det jag söker efter .
jag har fortfarande inte hittat det jag letar efter .
jag tycker att du behöver tänka på framtiden .
jag fick en bot på tjugo dollar för olovlig parkering .
jag såg på när de flådde en människa den dagen .
jag ser fram emot att få ditt brev .
jag ser fram emot sommarlovet .
jag är ledsen för hur jag betedde mig i går kväll .
jag är säker på att det skulle vara ett misstag att berätta för Tom .
jag är säker på att det vore ett misstag att berätta för Tom .
jag har gått och tänkte på det hela dagen .
jag har tänkt på det hela dagen .
jag har hört den franska versionen av den här låten .
på den tiden bodde han i huset ensam .
det spelar ingen roll vilket lag som vinner matchen .
klockan är nästan sju . vi måste gå till skolan .
att bo i en storstad har många fördelar .
malaria är en sjukdom som myggor bär på .
många träd tappar löven på vintern .
mor går till sjukhuset på morgonen .
en av tigrarna rymde från djurparken .
en av tigrarna rymde från zoot .
Julstjärnor är giftiga för katter och hundar .
hon lyckades inte övertala honom till att hålla tal .
hon var tvungen att dela sovrum med sin syster .
hon ser fram emot att få träffa honom igen .
någon måste vara här för barnen .
något kommer att hända . jag känner det på mig .
Förlåt , det hade jag fullständigt glömt bort .
tala högre så att alla kan höra dig .
schweizisk choklad smälter verkligen i munnen .
tack för chokladen . den var jättegod .
pojken som står vid dörren är min bror .
kyrkan står mitt i byn .
Regeringens politik misslyckades kapitalt .
Invånarna på ön är vänliga .
mannen erkände slutligen vad han hade gjort .
mannen erkände äntligen vad han hade gjort .
mannen erkände till slut vad han hade gjort .
mannen erkände till sist vad han hade gjort .
polisen tror att Tom förgiftade sig själv .
den stackars mannen blev äntligen en känd artist .
du har inget att vara arg över .
de här blommorna blommar tidigare än vad andra gör .
de är villiga att tala om problemet .
de har läst en intressant bok .
de är på god fot med sina grannar .
Tom och Mary har varit gifta i tre år .
Tom kunde knappt förstå vad Mary sade .
Tom förstår inte värdet av sparande .
Tom är den enda jag vet som kan göra det här .
Tom är den enda jag känner till som kan göra det här .
Tom är den enda jag vet om som kan göra det här .
Tom är för dum för att förstå dina skämt .
Tom tog ut en penna och började skriva .
Tom tog fram en penna och började skriva .
Tom gick in på sitt rum och stängde dörren .
två män med skidmasker gick in i banken .
var det dig jag hörde sjunga i duschen ?
vi blev väldigt besvikna över att höra nyheterna .
vi kommer inte att hinna , eller hur ?
vilken är din favoritsnabbmatsrestaurang ?
vad för slags amerikansk accent har Tom ?
vad skulle världen vara utan kvinnor ?
vad vill du bli när du blir stor ?
vilket år var det Berlinmuren föll ?
du har ingen aning om hur mycket det betyder för mig .
din högra strumpa är utochinvänd .
du måste stå i en kö för att köpa biljetten .
till att börja med borde du inte ha kommit hit .
Atomenergi kan användas för fredliga ändamål .
kom in . vi skulle precis sätta igång .
kom in . vi ska precis sätta i gång .
sa Tom något om det till dig ?
vill du inte höra min sida av historien ?
vill ni inte höra min sida av historien ?
vill du inte höra min syn på saken ?
vill ni inte höra min syn på saken ?
vill du inte höra min sida av saken ?
vill ni inte höra min sida av saken ?
vill du inte höra min version ?
han kunde inte förmå sig att skjuta hjorten .
han sover under dagarna och jobbar under nätterna .
hur fick du tag på en sådan stor summa pengar ?
hur vet jag om en tjej är intresserad av mig ?
hur lång tid tar det till stationen ?
hur många syskon har Tom ?
hur många dagar vill du vara i Boston ?
hur många dagar vill du tillbringa i Boston ?
hur många galaxer finns det i universum ?
jag är ekonomiskt oberoende av mina föräldrar .
jag såg på honom att han bara låtsades läsa .
jag tycker inte om honom , för han är slug som en räv .
jag tycker inte om sporter som tennis och golf .
jag vet inte vad som kommer att hända .
jag vill inte sjunga , för jag är tondöv .
jag fick schampo i ögonen och det svider .
jag hoppas att få se renar under min resa till Sverige .
jag vill bara vara din vän , ingenting mer .
jag tänker gå . jag bryr mig inte om du tänker göra det eller inte .
jag tänker åka . jag bryr mig inte om du tänker göra det eller inte .
jag spelade schack med Tom igår eftermiddag .
jag vill verkligen inte lämna barnen ensamma nu .
jag borde ha vetat bättre än att ringa honom .
jag tror jag aldrig har sett dig så full förut .
jag tycker att vi ska vänta en halvtimme till .
jag var i området , så jag tänkte komma förbi .
jag blev kidnappad när jag var tolv år gammal .
jag var inte medveten om att du mådde så dåligt .
jag åkte till Italien för andra gången 1980 .
jag skulle vilja betala med mitt kreditkort i stället .
jag vill att du går på mötet imorgon .
jag struntar hellre i skolan och spelar tv @-@ spel istället .
jag ska ta med min son till djurparken i eftermiddag .
det var du som föreslog att vi skulle se den filmen .
det är faktiskt mycket enklare än vad det ser ut .
det är oartigt att fråga hur mycket någon tjänar .
vänta en sekund . detta telefonsamtalet kan vara viktigt .
Kyoto är känt för sina helgedomar och tempel .
min bil är stor nog för fem personer .
ingen kunde förklara hur saken var gjord .
man har funnit olja under Nordsjön .
vid hemkomsten upptäckte jag inbrottet .
vår engelsklärare är både sträng och snäll .
snälla ge mig ett plåster och lite medicin .
hon blandar ofta ihop socker och salt .
hon betalade sju procents ränta på lånet .
medicinen var hennes sista utväg .
hon har inte varit i skolan på fem dagar .
en dag skulle jag vilja äga en segelbåt .
att simma över sjön tog nästan kol på mig .
djuret kämpade för att ta sig ut ur buren .
Kassören stoppade kundens varor i en påse .
den ekonomiska situationen är inte bra just nu .
polisen stängde Toms lemonadstånd .
Fången var bakom galler i två månader .
läraren tolkade meningen åt oss .
vädret ska bli bättre imorgon .
det finns ett akut behov av bloddonationer .
det fanns inga radioapparater i Japan på den tiden .
det finns en svensk ambassad i Washington D.C .
de hade inga skägg , inget hår och inga ögonbryn .
de gjorde aldrig det de sa att de skulle göra .
de övertalade mig att stanna ett tag till .
den här boken är för mig vad Bibeln är för dig .
det här monumentet restes i februari 1985 .
Tom kommer att stanna i tre dagar till .
Tom stannar i tre dagar till .
Tom är väldigt intresserad av grekisk mytologi .
Tom vill bara ha en muffins och en kopp kaffe .
Tom äter ofta äggröra till frukost .
Tom hällde upp lite mjölk i en skål till sina katter .
Tom sade att han tyckte att jag verkade imponerad .
Tom tror att Mary kan ha en ätstörning .
Tom kommer att bo hos oss ett par veckor .
Toms födelsedag var i förrgår .
vi har varit strömlösa i tre dagar nu .
hur stor procent av alla giftermål slutar med skilsmässa ?
vem bryr sig om Tom äter äggulor eller inte .
du får inte komma in här om du inte har ett pass .
du måste ha blandat ihop mig med någon annan .
du borde inte döma folk efter utseendet .
ett jobb är inte enbart ett sätt att försörja sig .
sa Tom hur länge Mary skulle vara i Boston ?
få saker ger oss så mycket nöje som musik .
han anmärker alltid på andra människor .
han spelade golf varje dag under semestern .
han lovade mig att komma förbi senast fem .
han lovade mig att titta förbi senast fem .
han säger alltid elaka saker om sin fru .
hur lång tid tog det honom att skriva den här romanen ?
hur lång tid tog det honom att skriva denna roman ?
hur många prenumeranter har den här tidskriften ?
jag är hungrig eftersom jag inte åt frukost .
jag minns inte exakt var jag la nycklarna .
jag kommer inte ihåg exakt var jag la nycklarna .
Jeg vet inte om han kommer att besöka oss nästa söndag .
jag har inte sett av honom på ett tag .
jag vet att Mary är vackrare än jag är .
jag kunde inte föreställa mig att jag skulle känna såhär för dig .
jag fick reda på det av en ren händelse .
jag trodde att Tom skulle sova över i Boston .
jag tog för givet att du skulle ansluta dig till oss .
jag åkte till Europa via USA .
jag önskar att jag hade lärt mig franska som barn .
jag undrar om det finns tillräckligt med mat åt alla .
jag vill helst inte äta samma mat i dag igen .
jag är säker på att jag kommer vinna tennismatchen .
jag ska arbeta under sportlovet .
jag letar efter någon att förälska mig i .
jag söker efter någon att förälska mig i .
Förlåt att jag har orsakat dig så mycket besvär .
jag har aldrig hört dig klaga på någonting .
vill du inte sjunga , behöver du inte det .
om du inte vill sjunga , behöver du inte det .
1891 blev Liliuokalani Hawaiis drottning .
i det avseendet håller jag fullständigt med dig .
det är tydligt att han stal pengar från kassaskåpet .
det är tydligt att han stal pengar ur kassaskåpet .
det här är inte min åsikt , bara min översättning !
mitt hus ligger i norra delen av staden .
mina föräldrar följde med till flygplatsen för att vinka av mig
Kärnvapen är ett hot mot hela mänskligheten .
kaniner är besläktade med bävrar och ekorrar .
hon valde ut en rosa skjorta för mig att prova .
hon sa att de var goda vänner till henne .
en del pojkar spelar tennis och andra spelar fotboll .
Tjuvar bröt sig in i mitt hus i går kväll .
Skådespelarens karriär räckte trettio år .
Porslinet ställdes ut i ett speciellt vitrinskåp .
fienden kastade in nya styrkor i slaget .
Vindruvorna är så sura att jag inte kan äta dem .
frågan var omöjlig för oss att besvara .
det röda paraplyt påminde henne om sin farmor .
det röda paraplyt påminde henne om sin mormor .
skolan ligger en halv mils väg från mitt hus .
Väggarna i det gamla huset var inte raka .
under soffan finns många dammråttor .
det finns många dammråttor under soffan .
det finns folk som läser böcker för att slå ihjäl tid .
det ligger en fjärrkontroll till tv:n under soffan .
de säger att han har varit död i två år .
denna salen tar 2000 personer .
det här är en tropisk storm . den är snart över .
Tom frågade om någon visste något om Mary .
Tom känner inte för att prata just nu .
Tom satte sig i förarsätet och körde iväg .
Tom har ett bankkonto på Caymanöarna .
Tom är definitivt inte på skämthumör idag .
Tom ljuger . jag gjorde inte det som han sa att jag gjorde .
Tom är den ende man som Mary någonsin har älskat .
Tom säger att han är villig att göra det gratis .
Tom verkar inte vilja sänka priset .
Toms mamma sa åt honom att klippa sig .
vi blir tvungna att skjuta upp matchen till nästa söndag .
vi ska mötas på stationen klockan nio .
vem tog hand om hunden medan du var borta ?
vem tog hand om hunden medan ni var borta ?
varför tror du att jag tänker på dig ?
Arbetsnarkomaner ser semesterdagar som slöseri med tid .
Arbetsnarkomaner ser semester som tidsslöseri .
du kan alltid räkna med honom i en nödsituation .
du har bara en chans att svara rätt .
du verkar gilla det här lika mycket som jag .
du borde inte gå ut i den här kylan .
din fråga hör inte till ämnet .
en vacker tjej med svart hår var i parken .
en vacker flicka med svart hår var i parken .
Enligt nyheterna blev han uppäten av hajar .
alla kommande möten kommer att hållas i detta rum .
en av stålets viktiga egenskaper är dess hållfasthet .
faktum är att han inte håller med mig .
så vitt jag vet håller de alltid sina löften .
det visade sig att han visste allt om mig .
vet du varför han skolkade idag ?
vet du anledningen till att han skolkade idag ?
lägg inte plånboken ovanpå elementet .
Ärligt talat , jag är inte särskilt imponerad av hans idée .
han bröt sitt löfte , vilket var ett stort misstag .
han visste inte vad han skulle göra med den överblivna maten .
han skadades allvarligt i trafikolyckan .
han klagar jämt på sin låga lön .
han söker desperat efter fler bevis .
han är inte alltid på kontoret på morgonen .
han var snäll nog att köra mig till sjukhuset .
han såg på kapplöpningen med sin kikare .
hur länge tänker du stanna här i Brasilien ?
hur många spel har du i din samling ?
jag kan inte fatta att jag pratar med dig om det här .
jag kan inte fatta att jag pratar med er om det här .
jag tvättade medan spädbarnet sov .
jag tror inte att ungen kom till Tokyo själv .
jag förstår inte vad du pratar om .
jag går till biblioteket två till tre gånger om veckan .
jag går till biblioteket två eller tre gånger i veckan .
jag går till biblioteket två till tre gånger per vecka .
jag blev tvungen att vänta i tjugo minuter på nästa bus .
jag behöver gå ner i vikt , så jag håller på med en diet .
jag vill tro att jag vet vad jag pratar om .
jag tycker att killar som kan spela piano är coola .
du borde nog berätta för Tom att du älskar honom .
i framtiden vill jag bli en TV @-@ presentatör .
jag var inte medveten om att du mådde så dåligt .
jag ska gå rakt på sak . du får sparken .
jag ska prata med Tom när han kommer hem .
jag ser fram emot att få träffa dig nästa söndag .
jag är trött på att alltid behöva göra allt arbete .
jag har lärt Tom att spela gitarr .
jag har beslutat mig för att svara på alla frågor offentligt .
om Tom hade sett någonting , skulle han ha sagt det till oss .
hade Tom sett någonting , skulle han ha sagt det till oss .
hade Tom sett något , skulle han ha sagt det till oss .
på den tiden var det få som kunde resa utomlands .
på den tiden kunde få människor resa utomlands .
det behöver inte innebära att du har rätt .
det är skönt att stiga upp tidigt .
ibland är det svårt att skilja rätt från fel .
det är ett för svårt problem för mig att lösa .
det kommer att ta några dagar att gå in de här skorna .
många företag gör reklam för sina produkter på tv .
min dröm är att leva fredfullt i byn .
snälla sänk volymen lite till .
Plutonium @-@ 239 har en halveringstid på 24 100 år .
hon steg på bussen och satte sig långt fram .
hon steg på bussen och tog plats långt fram .
hon valde skorna som matchar klänningen .
hon verkar vara förtjust med att prata om sig själv .
några är dyra medan andra är väldigt billiga .
Vissa gillar kaffe och andra gillar te .
Vissa tycker om kaffe och andra tycker om te .
Vissa människor gillar kaffe och andra människor gillar te .
äpplena han skickade mig var utsökta .
matchen kan ha skjutits upp till nästa vecka .
flickan var snäll och berättade vägen till museet .
ön är sex gånger Manhattans storlek .
Domaren dömde honom till ett års fängelse .
den andra delen av boken utspelar sig i England .
situationen är mycket värre än vi föreställt oss .
situationen är mycket värre än vi hade föreställt oss .
situationen är mycket värre än vad vi föreställt oss .
Stormen fick allvarliga följder för ekonomin .
läraren skrev någonting på svarta tavlan .
världens största djurpark finns i Berlin , Tyskland .
det går inte att förutsäga vad som kommer hända nästa år .
det var få elever kvar i klassrummet .
dessa fabriker förorenar miljön .
det här är det sötaste spädbarnet jag någonsin har sett .
Tom tillsatte några intressanta kryddor i stuvningen .
Tom och Mary åt upp hela tårtan själva .
Tom och Mary åt upp hela kakan själva .
Tom ägnade hela sitt liv åt att studera hajar .
Tom förstod inte att han gjorde ett misstag .
Tom har två sönder . bägge bor i Boston .
Tom tittade Mary djupt i ögonen och log .
Tom försöker skriva ett nytt blogginlägg varje dag .
Olyckligtvis släppte Tom ut katten ur säcken .
Olyckligtvis försade sig Tom .
Olyckligtvis avslöjade Tom hemligheten .
vi känner till legenden om Robin Hood .
hur dags går nästa tåg till Tokyo ?
vad händer om det blir ett strömavbrott nu ?
vilken föredrar du ? den här eller den där ?
medan du kör , borde du ha fokus på vägen .
kan du ta hand om våra husdjur medan vi är borta ?
kan ni ta hand om våra husdjur medan vi är borta ?
det går inte att förväxla honom med hans lillebror .
du ser trött ut , så du borde gå och lägga dig tidigt .
ni ser trötta ut , så ni borde gå och lägga er tidigt .
du kommer inte kunna övertala Tom att göra det där .
du är det vackraste flickan jag någonsin sett .
du är den enda person jag känner som kan hjälpa mig .
&quot; vill du lämna ett meddelande ? &quot; &quot; nej , tack &quot; .
en bra lärare måste vara tålmodig med sina elever .
en man som kan två språk är värd två män .
ett gräl uppstod om vad som man skulle göra med marken .
en 90 @-@ gradig vinkel kallas en rät vinkel .
Boston har vuxit i snabb takt de senaste tio åren .
Boston har vuxit snabbt de senaste tio åren .
Generellt sett lever kvinnor längre än män .
väck Tom och säg att frukosten är färdig .
gå och väck Tom och säg att frukosten är färdig .
han kom till New York för att söka jobb .
han bestämde sig för att en gång för alla sluta röka .
han beskrev olyckan i detalj .
han gör misstag varje gång han pratar engelska .
han vann första pris på schackturneringen .
hur många ingenjörer deltog i konferensen ?
jag visste inte hur jag skulle svara på hans fråga .
jag uppfattade inte riktigt namnet på den där designern .
jag avskyr kvinnor som säger att alla män är likadana .
jag måste gå och handla . jag är tillbaka om en timme .
jag tycker om att simma , men inte här .
jag såg en väldigt intressant dokumentär igår .
jag föreslår att vi tar det lite långsammare den här gången .
jag tror att vi har köpt allt som vi behöver .
jag tror att vi valde fel person för jobbet .
jag trodde du var van vid att bo i husvagn .
jag vill att du berättar allt som hände .
jag vill att du berättar allting som hände .
jag är riktigt trött . idag gick jag alldeles för mycket .
om du tänker döda mig så vill jag veta varför .
är det något särskilt som du vill ?
det ryktas att det finns gömda skatter här .
det var inte förrän igår jag fick nyheterna .
det var inte förrän i går som jag nåddes av nyheten .
det var inte förrän i går som jag nåddes av nyheterna .
min bror hjälper mig med läxorna ibland .
mitt hus ligger tio minuters gångväg från stationen .
hon kan inte bara tala engelska , utan också franska .
hon kunde inte hindra sin dotter från att gå ut .
hon målar varje dag , oavsett hur mycket hon har att göra .
hon är nyfiken på att få reda på vem det var som skickade blommorna .
någon måste ha tagit mitt paraply av misstag .
barnen åt chokladpudding till efterrätt .
kaffet var så varmt så jag inte kunde dricka det .
Patientens skador är inte livshotande .
de senaste medicinska framgångarna är anmärkningsvärda .
det finns inga matbutiker i närheten .
det finns inte så många synagogor i den här stan .
det finns ingen reguljär båttrafik till ön .
de säljer diverse varor på den affären .
de säljer diverse varor i den affären .
Tom och Mary tittade bekymrat på varandra .
Tom tvivlar inte på Marys förmåga att utföra jobbet .
Tom går på en promenad varje morgon med sin hund .
Tom fick mig att lova att inte säga någonting till dig .
Tom sa att han trodde att Mary kunde svetsa .
Tom ville att jag skulle spela schack med honom , så det gjorde jag .
två tredjedelar av eleverna kom till mötet .
vi har inte bestämt ännu vart vi ska åka imorgon .
vi använder ätpinnar istället för kniv och gaffel .
när det gäller tennis är hon överlägsen .
varför inte ansöka om jobbet som tolk ?
kvinnor känner att män ofta är väldigt komplicerade .
du behöver en bra utrustning för att klättra upp för det där berget .
du borde ha avvisat ett sådant orättvist förslag .
en tjuv bröt sig in i huset när vi var borta .
en gammal man vilade sig i skuggan av trädet .
förresten , hur många av er för dagbok ?
bli inte sårad . Tom är så där med alla .
för tusende gången : jag behöver inte din hjälp .
jag planerar att bo på hotell tills vidare .
han komponerade en begravningsmarsch till sin egen begravning .
han hörde illa och kunde inte gå .
han var tvungen att lämna staden , så han flyttade till Berlin .
han tänkte att det skulle vara vettigt att acceptera erbjudandet .
han översatte Homeros från grekiska till engelska .
han arbetar som lärare , men egentligen är han spion .
jag står inte ut med tanken på att förlora dig för evigt .
jag mår inte bra . snälla ge mig lite medicin .
jag förstår inte varför folk tror på spöken .
jag glömde stänga av tv:n före jag gick och lade mig .
jag fick ett brev som underrättade mig om hans ankomst .
jag tog för givet att du var på vår sida .
jag vill äta koreansk mat som inte är kryddstark .
jag fick veta att du kände till Toms telefonnummer .
du får ursäkta , men jag vill helst inte prata om det .
om du inte studerar mer så kommer du helt säkert att misslyckas .
det låg inte i hans natur att tala illa om andra .
inte förrän då fick han reda på sanningen .
det kanske var Tom som stal Marys halsband .
fler och fler studenter ansluter sig till protesterna .
min pappa insisterade på att vi skulle vänta på tåget .
det råder ingen tvekan om att hon älskar honom , men hon vill inte gifta sig med honom .
en för alla och alla för en , det är vårt motto .
du kanske rent av vet mer om det här än vad jag gör .
hon skämdes för sin obetänksamhet .
den där blonda tjejen med lockigt hår är från Sverige .
det var första gången någonsin jag körde bil .
Themsen är en flod som flyter genom London .
läkaren rådde min pappa att sluta röka .
hunden var upptagen med att gräva ner sitt ben i trädgården .
Utforskarna upptäckte ett skelett i grottan .
sista ansökningsdag är i övermorgon .
de två männen som satt på bänken var amerikaner .
vinden var så kraftig att fönstren skallrade .
det finns många amerikaner som kan tala japanska .
de har ännu inte fastlagt datumet för sitt bröllop .
de började sälja en ny typ av bil i Tokyo .
det här är den vackraste blomman i trädgården .
Tom bär alltid en karta och kompass i sin väska .
Tom och Mary tittar på teve i vardagsrummet .
Tom vet inte ens hur man startar en gräsklippare .
Tom körde av vägen när han väjde för en hund .
Tom tog av sig rocken och kastade den på golvet .
Tom brukade röka två paket cigaretter varje dag .
vi fick aldrig någon tydlig förklaring på mysteriet .
du då ? vill du också ha apelsinjuice ?
du då ? vill du också ha apelsinjos ?
vad får dig att tro att Tom gillar heavy metal ?
vad är skillnaden mellan sylt och marmelad ?
när jag blir stor ska jag gifta mig med Tom .
du hinner inte i tid till skolan .
du borde säga det till din mamma så snart som möjligt .
du vänjer dig snart vid din nya skola .
en tesked malen kanel är ungefär två gram .
Enligt tidningen begick han självmord .
allt som är för dumt för att sägas sjungs .
vet du inte att han gick bort för två år sedan ?
alla säger att han ser ut precis som sin far .
ursäkta , kan du sänka rösten lite ?
ungefär 9,4 % av jordens yta är täckt av skog .
han ådrog sig malaria när han bodde i djungeln .
han gick upp tidigt för att han skulle komma i tid till tåget .
han återvände hem efter att ha varit borta under tio månader .
han sade att han skulle hem nästkommande dag .
han försökte att göra sin fru lycklig , men han kunde inte .
han var intresserad av Orientens mysterium .
hur fick Tom Mary till att dansa med honom ?
hur många julkort skrev du förra året ?
jag dricker alltid två koppar kaffe varje morgon .
jag minns inte exakt vad jag ska göra .
jag visste inte att Tom inte har ett körkort .
jag har en vän vars far är en känd pianist .
jag höll i repet hårt så att jag inte skulle falla .
jag höll hårt i repet så att jag inte skulle falla .
jag sätter in tiotusen yen på banken varje månad .
jag vill ha en båt som kan ta mig långt härifrån .
jag vill äta något som jag bara kan äta här .
jag är inte säker på att det kommer att hända när som helst snart .
jag har försökt att lösa det här problemet i timmar .
trots att det regnade ställdes matchen inte in .
det gör ont att behöva säga det här , men det är sanningen .
det är inte nödvändigt för oss att närvara vid mötet .
det tog mig en halvtimme att lösa det här problemet .
det var inte nödvändigt att han skulle ta med ett paraply .
Seansdeltagare försöker få kontakt med de döda .
snälla låt mig få plocka upp din syster på stationen .
Skolor och vägar är tjänster som betalas för med skatter .
hon såg till att resenären hade mat och kläder .
hon höll just på att skära upp gurkor .
en del döva personer väljer att inte använda teckenspråk .
säg mig vad du äter , så ska jag säga dig vad du är .
Biskopen förbarmade sig över de förtvivlade immigranterna .
faktum är att hon läste inte ens brevet .
sjön hade frusit till , så vi gick över isen .
den gamla kvinnan gick upp för trappan med möda .
Offret låg med ansiktet ned i mattan .
det här skrivbordet som jag köpte igår är väldigt stort .
det här är den vackraste solnedgång jag någonsin sett .
i dag är morgondagen som vi oroade oss för i går .
i dag är morgondagen vi oroade oss för i går .
Tom frågade mig om jag verkligen trodde att jag kunde göra det
Tom kunde inte sova för han hade väldigt ont i huvudet .
Tom kunde inte sova för han hade en kraftig huvudvärk .
Tom ville inte skriva om det som hade hänt .
Tom tömde papperskorgen i förbränningsugnen .
Tom sade att han tyckte att jag verkade imponerad .
Tom satt tålmodigt i sin stol och väntade på Mary .
Tom ville bli teckenspråkstolk .
vi klev upp tidigt så att vi kunde se soluppgången .
vi steg upp tidigt så att vi kunde se soluppgången .
vi måste försöka att få in alla i huset .
ser du efter barnen medan jag är ute ?
i går köpte jag tio nya par ankelsockor .
du går inte upp lika tidigt som din syster , eller hur ?
du var med Tom natten han dog , eller hur ?
&quot; varför ska du inte åka ? &quot; &quot; för att jag inte vill &quot; .
&quot; varför ska du inte åka ? &quot; &quot; för jag vill inte &quot; .
Sömnbrist påverkade sångarens uppträdande .
alla äpplen som faller till marken äts upp av grisarna .
hur som helst , det kommer att vara en bra erfarenhet för dig .
känner du någon som var på det där skeppet som sjönk ?
hans försök med att simma över floden misslyckades .
han misslyckades med att försöka simma över floden .
han har setts som Japans svar på Picasso .
jag tänker skriva om våra parker och berg .
jag odlade tomater förra året och de smakade väldigt gott .
jag odlade tomater förra året och de var väldigt goda .
jag avskyr att ha med kräsna barn att göra .
jag behöver förstå vad denna mening betyder .
jag önskar bara att jag kunde vara så lycklig som du verkar .
jag trodde att Tom skulle tala bättre franska än Mary .
jag tog det för givet att du skulle följa med .
jag tänkte ringa honom , men jag kom på bättre tankar .
jag skulle aldrig ha gissat att Tom är från Boston .
det har tagit fyrtiosex år att bygga det här templet .
antingen talar vi kinesiska , eller så talar vi inte alls .
att förlora min dotter har berövat mig livsglädjen .
min mormor bor i Osaka .
min storebror lånade pengar av en kredithaj .
min storebror lånade pengar av en ockrare .
vår engelsklärare lägger vikt vid uttalet .
president Truman var tvungen att fatta ett svårt beslut .
president Truman var tvungen att ta ett svårt beslut .
hon hjälpte sin far med trädgårdsarbetet .
hon rörde om pulverkaffet och hällde i mjölk .
hon varnade barnen för att leka på gatan .
sluta gå som katten kring en het gröt och kom till saken .
den psykiatern har specialiserat sig på ätstörningar .
folkmassan demonstrerade för mänskliga rättigheter .
den officiella middagen ägde rum i Vita huset .
repet gick av medan vi besteg berget .
skolan är på gångavstånd från mitt hus .
Förhandlingarna ska ta upp problemet om miljöförorening .
det finns ännu några vilda folkstammar på den där ön .
Tom och hans bror klipper vanligtvis varandras hår .
Tom och hans bror klippte vanligtvis varandras hår .
Tom tycker inte om sättet hans mamma klipper hans hår på .
Tom har bestämt sig för att inte klippa sig förrän till våren .
Tom sa att han ville komma bort från stan ett tag .
Tom sade att han ville komma bort från staden ett tag .
Tom verkar ha hamnat i något slags koma .
ni verkade inte förstå vad Tom sa .
ni behöver inte förstå allt just nu .
du måste ta med dig ditt pass till banken .
du verkar ha förväxlat mig med min storebror .
du ska alltid skydda dina ögon från direkt solljus .
du jobbar för hårt . ta det lugnt en stund .
Zürich betraktas som en större finansiell knutpunkt .
en sexsiffrig inkomst är inte ovanligt för en läkare .
minns du när du vaknade i morse ?
han håller alltid fast vid att ha allting på sitt sätt .
han tappade kontrollen över bilen i kurvan .
jag antar att du jobbar på att rätta felen .
jag mår inte bra idag och föredrar att stanna hemma .
jag mår inte så bra . skulle du kunna ge mig lite medicin ?
jag tror inte att tv någonsin kommer att ersätta böcker .
jag hade en intressant konversation med min granne .
jag hatar när mina kläder luktar cigarettrök .
jag tror att vi köpt så gott som allt vi behöver .
jag tittade på en film på franska med engelska undertexter .
jag skulle vilja utbyta några ord med Tom i enrum .
jag skulle vilja tala ett slag med Tom mellan fyra ögon .
jag letar efter en man som ska bo här .
jag har skrivit ned alla siffror upp till trettioett .
det är svårt för en nybörjare att uppskatta vindsurfing .
deras kontor visade sig ha många kvinnor .
många unga i Japan äter bröd till frukost .
New York är en av de största städerna i världen .
ingen med namnet Tom Jackson har blivit anmäld som saknad .
hon bad mig att se efter hennes bebis medans hon var borta .
hon dukade av bordet efter middagen .
hon har studerat engelska sedan tioårsåldern .
hon pratar engelska som om det vore hennes modersmål .
tack för att du accepterade min vänförfrågan på Facebook .
namnet på de som dog har inte tillkännagetts .
de vill att vi ska tro att vi lever i en demokrati .
det här är kulan som läkaren tog ut från Tom .
det här är kulan som läkaren tog ut ur Tom .
detta är huset jag bodde i när jag var barn .
det här är den genväg som jag oftast tar till skolan .
det här är den genväg som jag brukar ta till skolan .
det här är genvägen jag brukar ta till skolan .
det här är den genväg till skolan som jag brukar ta .
detta är inte ett särskilt bra jobb , men det betalar räkningarna .
det är inte ett jättebra jobb , men det betalar räkningarna .
Tom lade inte märke till att Mary satt ensam .
Tom märkte inte att Mary satt ensam .
Tom sa att han skulle göra nästan vad som helst för Mary .
Tom såg festen som ett bra tillfälle att skapa nya kontakter .
vad är det för skillnad mellan en by och en stad ?
när han åker till Europa kommer han att besöka många museer .
Wikipedia är den bästa encyklopedin på nätet .
du kunde räkna till tio redan då du var två år gammal .
du pratar så fort att jag inte förstår ett ord av vad du säger .
du är den enda personen jag känner som inte äter kött .
ditt svar på frågan visade sig vara fel .
kan du säga mig hur man går till amerikanska ambassaden ?
vet du vilken gud det här templet är tillägnat ?
känns det bättre nu när du sovit en stund ?
bakterier kan bara ses med hjälp av ett mikroskop .
han övar på att spela gitarr tills sent på kvällen .
han skulle hellre dö än att gå upp tidigt varje morgon .
jag stannar här till i övermorgon .
jag fattar inte hur jag kunde tro att Tom skulle ändra på sig .
jag står inte ut med tanken på att förlora Tom som vän .
jag kan inte ta hennes plats som engelsklärare .
jag har precis varit på stationen för att vinka av min farbror .
jag har precis varit på stationen för att vinka av min morbror .
jag protesterade när kyparen försökte ta min tallrik .
jag brukade simma i havet när jag var ett barn .
jag ska ta körkort när jag blir arton .
jag skulle kunna förklara det för dig , men din hjärna skulle explodera .
jag skjuter upp min resa till Skottland tills det blir varmare .
om inte den där gitarren vore så dyr , så skulle jag kunna köpa den .
om du är upptagen nu kan jag ringa tillbaka till dig senare .
är det någon här som känner någon i Australien ?
det gör ont att behöva säga det här , men det är sanningen .
det tar oss fem minuter att gå igenom tunneln .
det tog honom tre månader att lära sig cykla .
det var hans bil , och inte min , som gick sönder i går .
det var snudd på otänkbart att pojken skulle stjäla .
det var snällt av dig att hjälpa mig med läxan .
det skulle inte förvåna mig om Tom och Mary gifte sig .
Oavsätt hur mycket hon äter , så går hon aldrig upp i vikt .
oavsett vad som händer kommer jag aldrig att ändra mig .
smärta är något vi alla måste lära oss att hantera .
folk ändras . det finns inte mycket du kan göra åt det .
var snäll och vänta en stund medan jag gör klart ditt kvitto .
Skolbarn är förkylda dubbelt så ofta som vuxna .
hon har sönder något varje gång hon städar rummet .
hon höll honom som gorillamammor håller sina ungar .
Förenta nationerna är en internationell organisation .
regeringen föll efter en omröstning i riksdagen .
Liftarna var närapå förfrusna när de hittades .
modern och dottern representerade två generationer .
den blyga pojken var ytterst generad i hennes närvaro .
läraren underströk vikten av att föra anteckningar .
problemet är att vi inte har någonstans att vara ikväll .
det finns runt tretusen moskéer i Istanbul .
det var en vacker flicka med svart hår i parken .
det var en vacker tjej med svart hår i parken .
Tom slumrade till , sittandes i solen på sin veranda .
Tom hade aldrig sett en älg förrän han flyttade till Alaska .
vad ska du göra under sommarlovet ?
vad ska du göra på sommarlovet ?
när han kom tillbaka hem , sov barnen redan .
vem blir den nästa presidenten av USA ?
du måste förstå problemets omfattning .
ett slukhål har bildats mitt i motorvägen .
alla vägar som leder in till staden är fulla av bilar .
vet du varför vårrullar kallas för vårrullar ?
vet ni varför vårrullar kallas för vårrullar ?
vet du varför vårrullar kallas vårrullar ?
vet ni varför vårrullar kallas vårrullar ?
vet du varför vårrullar heter vårrullar ?
vet ni varför vårrullar heter vårrullar ?
engelska talas i många länder runt om i världen .
fastän det låter märkligt är det sant det hon sade .
Gymnaster är bland de vigaste av alla idrottare .
han klagar på det ena och det andra hela tiden .
han bestämde sig inte för att bli författare förrän han var trettio .
vad sägs om glass och chokladsås till efterrätt ?
jag bestämde mig för att jag inte ville ha mer med Tom att göra .
jag har en lång lista saker jag inte borde göra
jag hoppas att något bra händer innan dagen är över .
jag lånade honom lite pengar , men han har inte betalat tillbaka dem än .
jag bodde en vecka i Berlin hos en tysk familj .
om jag visste hennes namn och adress kunde jag skriva till henne .
om du inte vill säga någonting , behöver du inte det .
vill du inte säga någonting , behöver du inte det .
om ni inte vill säga någonting , behöver ni inte det .
visst är han ung , men han är mycket pålitlig .
det luktar som om någon har rökt här inne .
det var mycket svårare än jag hade förväntat mig .
det var inte så lätt som vi trodde att det skulle vara .
var god fyll i enkäten och skicka in den till oss .
Sedd från flygplanet ser ön väldigt vacker ut .
han ska övertala sin far att köpa en ny bil .
polisen häktade ett flertal misstänkta för förhör .
läraren demonstrerade idén med ett experiment .
du behöver inte vara rädd . han kommer inte att göra dig illa .
det fanns bara ett fall av vattenkoppor på skolan .
Tom gav upp sin dröm om att bli oceanograf .
Tom gav upp sin dröm om att bli djuphavsforskare .
Tom förväntade sig inte riktigt att Mary skulle svara på hans fråga .
Tom missade chansen att åka till Boston med Mary .
Tom låtsades inte förstå vad Mary sa .
Tom tog av sig sina kläder och gick in i duschen .
Toms hus är ungefär tre kilometer härifrån .
Toms hus ligger ungefär tre kilometer härifrån .
vad är skillnaden mellan kantonesiska och mandarin ?
när jag kom hem , upptäckte jag att jag hade tappat bort min plånbok .
varför provade du inte klänningen innan du köpte den ?
du behöver inte säga någonting du inte vill säga .
i det här skedet behöver ni inte förstå allt .
har du lite bröd ? jag ska mata duvorna .
han har spelat schack sedan han gick på high school .
han är stolt över att ha tagit examen vid Tokyo Universitet .
hur många olika pjäser är det i japanskt schack ?
jag lärde mig att cykla när jag var sex år gammal .
det kan hända att jag är hemma i kväll , men jag är inte säker än .
jag undrar om hon kommer ihåg mig efter alla dessa år .
jag ska gå och hämta lite kaffe . vill du ha en kopp ?
om du inte vill hålla tal , behöver du inte det .
vill du inte hålla tal , behöver du inte det .
om du inte vill dit , så åker vi inte dit .
är det något särskilt som du vill ha att äta ?
min far har slutat röka för sin hälsas skull .
Vissa studenter kommer inte att komma tillbaka nästa termin .
några studenter kommer inte att komma tillbaka nästa termin .
Tornet är trehundratjugoen meter högt .
det finns inte plats här inne för både Tom och Mary .
de överlevde trots att byggnaden förstördes .
Tom är vänsterhänt , men han skriver med höger hand .
vi kommer troligen inte att göra det igen på ett tag .
vi vill veta hur mycket det här projektet kommer att kosta oss .
det är inte tillåtet för kvinnor att köra bil i Saudiarabien .
du borde läsa en sådan bok som han läser just nu .
en liter mjölk innehåller ungefär trettio gram protein .
Enligt tv @-@ nyheterna har det skett en flygkrasch i Indien .
alla hästar är djur , men inte alla djur är hästar .
Barnaga är fortfarande tillåtet i många länder .
vill du gifta dig först eller skaffa barn först ?
har alla i Sverige blont hår och blå ögon ?
Läs inte vad som är i brevet . bara ge det till Tom .
Frukter och grönsaker är en väsentlig del av en balanserad kost .
har du någonsin fått höra vad som faktiskt hände den dagen ?
han har sålt sin bil , så han tar tåget till kontoret .
han har vanan att läsa tidningar under måltider .
han har bott på det där hotellet de fem senaste dagarna .
jag kan inte stänga av duschen . kan du kolla det åt mig ?
jag lyckas inte stänga duschen . kan du kolla på det åt mig ?
jag har varit bekant med henne i över 20 år .
jag vet att du har viktigare saker att tänka på .
jag vet att ni har viktigare saker att tänka på .
jag söker ett läppstift som passar med det här nagellacket .
är det något särskilt som du vill höra ?
det är kanske ingen bra idé att äta medan du springer .
det är upp till dig att bestämma om vi skall gå eller inte .
John F. Fitzgerald valdes till borgmästare i Boston år 1906 .
min engelsklärare rekommenderade mig att läsa dessa böcker .
min engelsklärare rekommenderade mig att läsa de här böckerna .
folk säger ofta att japanska är ett svårt språk .
du kanske kan föreslå något vi kan göra imorgon .
hon tog på sig sin systers jeans och tittade i spegeln .
hon tog på sig sin systers jeans och såg sig i spegeln .
köpcentret var fullproppat med semestershoppare .
Diktatorn hade den absoluta lojaliteten av alla hans medhjälpare .
Diktatorn hade alla sina medhjälpares fulla lojalitet .
ju mer du lär känna henne , desto mer kommer du att gilla henne .
tröjan Tom hade på sig idag hade hans mamma gjort .
det finns viktiga frågor som måste bli besvarade .
det står nu tre bilar parkerade framför vårt hus .
de skymtade mannen genom folkmassan .
Tom sa alltid att han ville lära sig spela mahjong .
Tom kan inte tala franska . Mary kan inte heller tala franska .
Tom spenderade hela dagen med att designa en hemsida åt en ny kund .
Tom vaknade när han hörde någon knacka på dörren .
vi väntar oss många besökare till ceremonin .
vad är den bekvämaste vägen till Tokyo station ?
vilken är den bekvämaste vägen till Tokyo station ?
du har köpt fler frimärken än vad som är nödvändigt .
du borde koncentrera dig på vägen när du kör .
du var den vackraste kvinnan på festen ikväll .
du var den vackraste kvinnan på festen i kväll .
&quot; vad tänker du på ? &quot; &quot; jag tänker på dig &quot; .
som 90 @-@ åring lever Toms farmor fortfarande ett mycket aktivt liv .
både pojkar och flickor borde studera hemkunskap .
Gazpacho är en kall tomat- och grönsakssoppa från Spanien .
jag kunde inte ta mig utanför stadion på grund av folkmassan .
jag trodde aldrig att det skulle vara såhär svårt att skapa en iPad @-@ app .
om du pratar för snabbt , kommer jag inte att förstå .
är det något särskilt som du vill ha att dricka ?
är det något särskilt som du vill titta på ?
det är omöjligt att veta vad som kommer att hända i framtiden .
det var mörkt , så Tom hade problem med att läsa gatuskylten .
det erbjudandet låter för bra för att vara sant . vad är haken ?
presidenten ignorerade demonstranterna utanför sitt kontor .
de serverade inte Tom någon alkohol eftersom han var underårig .
det här är huset som jag bodde i när jag var liten .
det här är huset jag bodde i när jag var liten .
Tom låtsades inte höra Mary ropa hans namn .
Tom vaknade när han hörde någon knacka på dörren .
Toms hund lämnade leriga tassavtryck över hela hans nya matta .
vi har large , medium och small . vilken storlek vill du ha ?
vi har large , medium och small . vilken storlek vill ni ha ?
ska vi inte pausa en stund och dricka lite kaffe ?
när det regnar så här får vi aldrig en chans att gå !
alla skolungdomar går för halv priset under jullovet .
är du säker på att du inte vill stanna ett par dagar ?
kastanjer måste kokas i minst femton minuter .
barn vill höra samma historia om och om igen .
Cuzco är en av de intressantaste platserna i världen .
Etniska minoriteter kämpar mot fördomar och fattigdom .
han gick långsamt så att barnen skulle kunna klara av att följa efter .
jag har fortfarande kvar fotot jag tog på dig för 10 år sedan .
vi råkar ha två exemplar av &quot; Räddaren i nöden &quot; .
det är väldigt svårt att säga vilket land en person kommer ifrån .
det var aldrig svårt för oss att hitta något att prata om .
det var en av mitt livs mest makalösa upplevelser .
det vore bättre om du inte åt innan du gick till sängs .
föräldrar är ansvariga för sina barns säkerhet .
förr trodde man att bara människor kunde använda språk .
en del människor läser tidningen medan de ser på tv .
Premiärministern kommer att hålla en presskonferens imorgon .
Frihetsgudinnan är symbolen för USA .
pojken var så trött att han inte kunde ta ett steg till .
Nyhetsförmedlaren betonar matkrisen för mycket .
den förra hyresgästen skötte lägenheten utmärkt .
det här formuläret ser rätt komplicerat ut . hjälp mig att fylla i det .
det här är just den ordbok jag har letat efter .
det är just den här ordboken som jag har letat efter .
Tom och Mary gifte sig i oktober på en tropisk strand .
Tom visste inte att Marys hus var så nära Johns .
Tom säger att han inte har lust att dricka öl i kväll .
Tom var den ende som inte kunde franska .
vi kan inte bevisa att Tom ljuger , men vi är ganska säkra på att han gör det .
vad har det blivit av boken jag lade här för några minuter sedan ?
du kan komma och se mig närhelst det passar dig .
du behöver inte säga någonting om du inte känner för det .
ni behöver inte säga någonting om ni inte känner för det .
du behöver inte säga något om du inte känner för det .
ni behöver inte säga något om ni inte känner för det .
du behöver inte säga någonting om du inte har lust .
du behöver inte säga någonting om du inte har lust med det .
ni måste inte säga någonting om ni inte har lust .
en förbipasserande bil körde i en vattenpöl och stänkte ned hela mig .
kan du hjälpa mig att översätta dessa meningar till kinesiska ?
minns du första gången vi åkte till Boston tillsammans ?
han må vara ung , men han är verkligen en tillförlitlig person .
jag hade pluggat engelska i två timmar när han kom in .
jag har en vän vars far är kapten på ett stort skepp .
jag bodde i Tokyo för några år sedan , men nu bor jag i Kyoto .
jag minns att jag var på ett skepp när jag var bara fem år gammal .
jag trodde att Tom skulle plantera de där blommorna nära eken .
jag fick veta att du kunde lära mig hur man slipar en kniv .
om en dörrvakt bär ditt bagage , glöm inte att ge honom dricks .
det här är första gången jag skriver ett brev på spanska .
det är dags att inse att det är omöjligt . vi kommer aldrig att klara det .
oavsett hur snabbt du kör hinner du inte dit i tid .
vår lärare försökte att använda en ny metod för att lära ut engelska .
detta är ett litet steg för en människa men ett jättekliv för mänskligheten .
ett litet steg för en människa , ett stort steg för mänskligheten .
så fort som tjejen såg sin mamma så började hon att böla .
Korsningen där olyckan inträffade ligger här i närheten .
ön är täckt av is och snö under vintern .
polisen övertalade förbrytaren att lämna ifrån sig sitt vapen .
det går tre elever med samma namn i den klassen .
det finns ingenting på jorden som inte påverkas av solen .
det står en man med en pistol i handen i dörren .
det står en man med en pistol i handen vid dörren .
här är en mening , med stavelseantalet , som i en haiku .
Tom råkade skära sig i handen när han skivade morötter .
Tom äter yoghurt med hackad mandel på till frukost .
Tom är inte en lat pojke . i själva verket arbetar han hårt .
Tom rullade ihop affischen och stoppade in den i ett papprör .
Tom räddade Mary &apos; s liv genom att utföra Heimlichmanövern .
byggdes denna mur för att hålla människor ute eller för att hålla dem inne ?
byggdes denna mur för att hålla människor ute eller inne ?
byggdes den här muren för att hålla folk ute eller för att hålla dem inne ?
vi måste bränna alla de här grejerna innan polisen kommer .
en bra mening är inte nödvändigtvis en bra exempelmening .
en bra mening behöver inte vara en bra exempelmening .
alkohol löser inga problem , men det gör inte mjölk heller .
Jämför de båda noggrant , så ska du se skillnaden .
till och med under arbetstid ger jag i lönndom efter för mitt internetberoende .
han lovade mig att vara mer försiktig i framtiden .
hur visste du att jag skulle ställa den frågan till dig ?
hur många barn vill du ha när du gifter dig ?
hur gammal var du när du slutade tro på tomten ?
hur gamla var ni när ni slutade tro på tomten ?
hur gammal var du när du slutade tro på jultomten ?
hur gamla var ni när ni slutade tro på jultomten ?
jag är trött eftersom jag var tvungen att plugga inför ett prov igår natt .
jag får känslan av att ingen här berättar sanningen för oss .
jag hoppas att Tom stannar i Boston åtminstone tre dagar till .
jag visste att det skulle bli svårt att övertala Tom att hjälpa oss .
jag vill veta varför du inte gjorde det du sa att du skulle göra .
om du inte har något snällt att säga , säg ingenting alls .
om du någonsin kommer till Boston , är du välkommen att bo hos oss .
istället för att åka till Australien vill jag åka till Nya Zeeland
säg till henne att du gillar henne . var inte rädd . hon kommer inte att bita dig .
Avståndet från mitt hus till ert hus är två kilometer .
dimman var så tjock att jag inte kunde se vart jag var påväg .
det här kommer att bli den varmaste sommaren på trettiosex år .
Toms mamma sa alltid till honom att han borde äta mer grönsaker .
vad är skillnaden mellan amerikansk och brittisk engelska ?
skulle du kunna vakta den här väskan åt mig en liten stund ?
efter att ha misslyckats två gånger i går vill han inte försöka igen .
jag minns inte exakt hur gammal jag var när jag träffade Tom för första gången .
jag kommer inte ihåg hur gammal jag var när jag träffade Tom för första gången .
jag minns inte hur gammal jag var när jag för första gången träffade Tom .
jag kommer inte ihåg hur gammal jag var när jag för första gången träffade Tom .
jag får svår prestationsångest före jag ska hålla ett tal .
jag har en katt och en hund . katten är svart och hunden är vit .
jag tror att det är osannolikt att Tom kommer till festen själv .
det var nån som sa att Tom hade varit med om en trafikolycka .
på tal om tv , vilket är ditt favoritprogram nuförtiden ?
Britterna trodde att amerikanerna överträdde deras lag .
Britterna tyckte att amerikanerna överträdde deras lag .
Rockkonserten ställdes in , för sångaren blev sjuk .
de sa till Tom att han måste skriva under ett sekretessavtal .
det här är den kallaste vintern som vi har haft på trettio år .
Tom räddade hunden ifrån att bli uppäten av de hungriga soldaterna .
Tom sa att han brukade åka till Australien tre gånger om året .
vi måste lasta ur den här lastbilen innan det börjar regna .
när jag ser tillbaka på den där tiden verkar allt som en dröm .
igår var han väldigt sjuk men idag mår han mycket bättre .
hans utställning på stadsmuséet tilltalade mig inte alls .
hur många självmord tror du att det sker varje år i Japan ?
är det etiskt att ge honom intervjufrågorna i förväg ?
det var en så kraftfull explosion att taket flög av .
det var inte så svårt att göra som jag trodde det skulle vara .
min morfar dog för 10 år sedan .
eftersom jag hade träffat honom en gång innan , kände jag genast igen honom .
Trädgårdsmästaren planterade en ros mitt i trädgården .
det fanns mycket som vi helt enkelt inte hade tid att göra .
det här företaget använder billig arbetskraft för att öka sina vinstmarginaler .
det här var första gången någonsin Tom hade sett ett skrotbilsrally .
Tom klipper sig oftast bara två eller tre gånger om året .
Tom var den ende som inte lämnade in hemuppgifterna i tid .
Toms fru gillar inte när han röker i vardagsrummet .
vi förknippar namnet Darwin med evolutionsteorin .
Burj Khalifa är för närvarande världens högsta skyskrapa .
Burj Khalifa är för närvarande den högsta skyskrapan i världen .
Skyll inte på mig . jag har ingenting att göra med den där videon .
hennes frågor visar att hon är väl insatt i ämnet .
jag har en katt och en hund . katten är svart och hunden är vit .
jag hörde att en sydamerikansk campare blev uppäten av en anakonda .
om vädret är bra i morgon , går vi till floden och badar .
om vädret är bra i morgon , går vi till floden och simmar .
mina favoritämnen i gymnasiet var geometri och historia .
mina favoritämnen på gymnasiet var geometri och historia .
hon tittade på några klänningar och valde ut den dyraste .
hon säger att hon inte dejtar någon just nu , men jag tror inte på henne .
problemet är att pojken aldrig gör vad han blir tillsagd att göra .
till hela stadens förvåning , arresterades borgmästaren .
Tom kan inte sitta i bilen längre än tio minuter innan han blir åksjuk .
vi måste ta reda på om vi har tillräckligt med pengar för att göra det .
vi hinner förmodligen inte göra klart det idag .
du borde inte säga såna saker när barn är i närheten .
en färsk undersökning visar att antalet rökare minskar .
jag vill bara kunna besöka mina barn när jag så önskar .
jag vill bara kunna besöka mina barn när jag vill .
jag är rädd att jag inte kan göra mig förstådd på franska .
det kostade mig tiotusen yen att få min tv @-@ apparat reparerad .
att mingla med folk på fester kan vara förskräckande för blyga människor .
när man har fått in en dålig vana , så är det inte enkelt att bli av med den .
Öns ekonomi är beroende av fiskeindustrin .
Varorna som beställdes från England förra månaden har inte anlänt än .
här är en mening , med stavelseantalet , som i en haiku .
Tom låg vaken länge och tänkte på vad han skulle göra .
Tom låg vaken länge och tänkte på vad han borde göra .
Tom satt tre decennier i fängelse för ett brott han inte begick .
jag fick veta att det var svårt för henne att lösa det problemet .
jag försöker komma på varför någon skulle göra något sådant .
jag försöker komma på varför någon skulle göra någonting sådant .
jag försöker komma på varför någon skulle få för sig att göra något sådant .
jag försöker komma på varför någon skulle få för sig att göra någonting sådant .
Förlåt att jag ringer så sent . jag ville bara höra din röst .
att äta en klyfta vitlök varje dag , är det nyttigt för dig ?
är det bra för hälsan att äta en vitlöksklyfta om dagen ?
lista de fem bästa sakerna du gillar att göra när du inte jobbar .
Schweiz är ett väldigt vackert land och är mycket värt att besöka .
bron mellan Danmark och Sverige är nästan åtta kilometer lång .
Tom rådde Mary att inte tro på allt hon läser på webben .
Tom tillrådde Mary att inte tro på allt hon läser på webben .
Tom och Mary vaknade tidigt för att se årets första soluppgång .
Tom tittade ut genom fönstret på skeppet som kom in i hamnen .
Tom sa att han trodde att Mary fortfarande bodde hos sina föräldrar .
Tom tog av sig rocken eftersom det var för varmt för att ha den på sig .
Toms nya skjorta krympte i tvätten så nu passar den inte .
medan han pratade hördes ljudet av ett skott som avlossades .
medan han pratade hördes ett skott avlossas .
en förbipasserande filmade polisens våld med sin mobiltelefon .
kan du snälla säga hur lång du är och hur mycket du väger ?
elföretag försöker minska sin kolförbrukning .
jag hade hans namn på tungan , men jag kunde inte komma ihåg det .
jag sa till henne en gång för alla att jag inte skulle gå och handla med henne .
om du inte håller dina löften , kommer folk inte att ta dig på allvar .
på den tiden var Amerika inte självständigt från Storbritannien .
hon sa själv att hon inte skulle bli kär i någon igen .
det här ser ut att kunna vara vapnet som användes för att döda Tom .
Tom visade mig dikterna han skrev när han var tonåring .
två vuxenbiljetter och tre barnbiljetter till London , tack !
du kan se den stora utställningen på köpcentret vilken tid som helst .
en man som inte spenderar tid med sin familj kan inte vara en riktig man .
jag kan inte komma på någon bra ursäkt till varför jag är sen till tandläkaren .
jag sov inte bra i natt , så jag har inte så mycket energi i dag .
om du skulle prata mindre och lyssna mer , skulle du kanske lära dig någonting .
om du pratade mindre och lyssnade mer , skulle du kanske lära dig någonting .
hon höll kattungen som en gorillamamma skulle hålla sin egen unge .
skeppet genomsöktes noggrant , men inga illegala droger hittades .
det flyger en reklamballong ovanför köpcentret .
Tom satt vid poolen och drack rödvin och åt dyr ost .
&quot; hur lyckades ni bryta er in utan dyrk ? &quot; &quot; Toalettfönstret var öppet &quot; .
han har skaffat sig vanan att stoppa händerna i fickorna .
jag behöver inte gå till doktorn längre . jag mår mycket bättre .
jag träffade någon häromdagen som jag tror att jag skulle kunna bli kär i .
jag misstänkte att han ljög , men det kom inte som en överraskning .
jag undrade bara om du har lyckats hitta någonstans att bo .
det tog mig mer än två timmar att översätta några sidor i engelska .
det tog mig mer än två timmar att översätta några sidor engelska .
jag är på ett gräsligt humör i dag för jag har inte tillräckligt med pengar .
stanna gärna kvar efter konserten . vi kommer att skriva autografer .
hon hade precis börjat läsa boken när någon knackade på dörren .
Schweiz är beläget mellan Frankrike , Italien , Österrike och Tyskland .
jag har massor av begagnade böcker till salu , allt till överkomliga priser .
hon köper allt hon vill ha utan att bry sig om priset .
läkarna säger att det var ett mirakel att Tom överlevde natten .
antalet européer som besöker Thailand varje år , är mycket stort .
de exporterar mycket frukt såsom apelsiner , grapefrukter och citroner .
Tom vill inte bli läkare , trots att han är väldigt på naturvetenskap .
Tom ligger i koma och läkarna är inte säkra på om han kommer att överleva .
han uppskattar att det nya huset kommer kosta ungefär trettio miljoner yen .
jag kan inte komma på något annat sätt att få honom att acceptera vårt förslag .
Troligt är att inget språk fullständigt saknar lånord .
Mary satte några blommor i vasen och ställde sedan vasen på bordet .
Invånarna i staden är beroende av floden för att få dricksvatten .
Tänk på hur mycket värre det hade kunnat vara om Tom inte hade varit där .
det finns inget annat att göra än att vänta på att platserna blir lediga .
kan du förklara skillnaden mellan svart te och grönt te för mig ?
Etniska minoriteter kämpar mot fördomar , fattigdom och förtryck .
Långdistanslöpare är i allmänhet ovigare än kortdistanslöpare .
jag föreslår honom till ordförande oavsett om du är för det eller inte .
om hon bara hade vetat att jag var i Tokyo , skulle hon ha hälsat på mig .
företaget jag arbetade för höll på att skära ner . Olyckligtvis förlorade jag jobbet .
Tom tar en snabb joggingtur runt kvarteret varje morgon innan frukost .
hela dagen var min pappa på dåligt humör för att han tappat bort sin plånbok .
till följd av konstant hunger och utmattning dog hunden till slut .
det förvånar mig att Tom inte ens kan sjunga en enda sång på Franska .
vänlighet är det språk som de döva kan höra och de blinda kan se .
de flesta barn slutar att kissa i sängen vid sju eller åtta års ålder .
hon rådde honom att gå till sjukhuset , men han lydde inte hennes råd .
Tom frågade Mary några mycket personliga frågor som hon vägrade svara på .
Tom är levande bevis på att man inte behöver förstånd för att bli framgångsrik .
Olyckligtvis var min granne med om en trafikolycka och hamnade i koma .
före andra världskriget gick gränsen mellan Finland och Sovjetunionen nära Leningrad .
han växte upp i USA , men hans modersmål är japanska .
de två länderna hade stridit tillsammans som allierade under andra världskriget .
som pojke brukade jag ligga på gräset och titta på de vita molnen .
jag visste att jag var tvungen att berätta sanningen för honom , men jag kunde inte förmå mig till det .
hon tilläts att gå till discot , på villkor att hon var tillbaka vid tio .
för att bli en bra översättare så tror jag att Tom behöver finslipa sina kunskaper lite till .
Tom raderade av misstag alla filer på en av sina externa hårddiskar .
Toms farfar och Marys farfar slogs tillsammans i andra världskriget .
Toms farfar och Marys morfar slogs tillsammans i andra världskriget .
Toms morfar och Marys farfar slogs tillsammans i andra världskriget .
Toms morfar och Marys morfar slogs tillsammans i andra världskriget .
han betonade att tiotusentals människor skulle komma till konserten .
min far är stolt över det faktum att han aldrig varit i en trafikolycka .
jag har fyra datorer , men två av dem är så gamla att jag inte använder dem längre .
tycker du fortfarande att jag är den som du vill tillbringa resten av ditt liv med ?
efter att ha gått ur duschen , så torkade Tom bort dimman från spegeln och rakade sig .
jag tycker att vi ska göra som Tom föreslår , om inte någon annan har ett bättre förslag .
min farfar firar sin åttioåttonde födelsedag i morgon .
min morfar firar sin sextionde födelsedag i morgon .
hon höll kattungen på samma sätt som en gorillamamma skulle hålla sin egen unge .
vad har du för bevis på att det var Tom som stal din mors halsband ?
på grund av den dåliga skörden har vetepriset gått upp de senaste sex månaderna .
tror du att Tom faktiskt hade tänkt dricka hela vinflaskan själv ?
andra forskare diskuterar hans teori om dinosauriernas försvinnande .
sedan jag återhämtade mig från min allvarliga sjukdom ter sig hela skapelsen vacker för mig .
Barcelona är huvudstaden i Katalonien , och det är den näststörsta staden i Spanien .
du pratar lite för snabbt för mig . skulle du kunna prata lite långsammare ?
&quot; snön är vacker , eller hur ? &quot; &quot; ja , men Mary , du är ännu vackrare &quot; .
jag hade aldrig kunnat gissa att Tom och Mary skulle bli kära i varandra .
vi har inte mycket pengar , men vi har tillräckligt för att köpa det vi absolut behöver .
trots att jag har läst engelska 6 år i skolan talar jag det inte bra .
har du en minut ? jag skulle vilja diskutera någonting som är angeläget för oss båda .
Studier har visat att det genomsnittliga tangentbordet har mera bakterier än en toalettstol .
när jag besökte deras lägenhet , var paret mitt i ett gräl .
när jag gick i skolan blev vänsterhänta barn tvingade att skriva med höger hand .
min favoritsmoothie är en som är gjord på grönt te , frysta hallon och blåbär .
alla blev mycket förvånade över avslöjandet att slavflickan i själva verket var en prinsessa .
jag hörde att Tom hade smugglat droger till Amerika i flera år innan han åkte fast .
i medicinsk forskning är ett av de största problemen att ta reda på orsaken till sjukdomen .
om inte människan tar hand om miljön kanske miljön eliminerar mänskligheten .
en grundlig kännedom om datorsystem och programmeringsspråk är en väsentlig del av Toms arbete .
Tom bar nackkrage i flera månader efter att ha fått en pisksnärtskada i en bilolycka .
en kraftig man med ett mörkt utseende ryckte Marys handväska och försvann in i folkmassan .
föräldrar bokstaverar ofta ord och meningar som de inte vill att deras unga barn ska förstå .
popcorn är väldigt billigt , jämfört med många andra snacks . det är även oftast hälsosammare .
min far , farfar , farfars far och farfars farfar hade alla samma namn som jag .
på inrådan av sina astronomer bestämde sig Alexander den store för att inte attackera Egypten och for till Indien istället .
alla har rätt till sin egen åsikt . men ibland är det bättre att hålla den för sig själv .
Tom försökte sälja sin gamla videobandspelare istället för att slänga den , men ingen köpte den , så det slutade med att han slängde den .
Tom sa att han inte var intresserad av Mary , men det verkade som att han alltid tittade åt den del av rummet som hon var i .
när jag läste till jurist sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på .
när jag läste till advokat sa mina lärare åt mig att aldrig ställa en fråga som jag inte visste svaret på .
din engelska är grammatiskt riktig , men ibland låter det du säger bara inte som något en modersmålstalare skulle säga .
din engelska är grammatikalisk , men ibland låter det som du säger bara inte som någonting som en modersmålstalare skulle säga .
ett sätt att minska antalet fel i Tatoebas korpus skulle vara att uppmuntra människor att endast översätta till sina modersmål .
ett sätt att minska antalet fel i Tatoebas korpus vore att uppmuntra människor att endast översätta till sina modersmål .
ett sätt att minska antalet fel i Tatoebas korpus vore att uppmuntra folk att endast översätta till sina modersmål .
om du tar med ett barn ut och pekar på månen , så tittar barnet på månen . gör du samma sak med en hund så tittar den på ditt finger .
