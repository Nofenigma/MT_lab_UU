ge mig en sekund .
det är ett av mina favoritord .
han gillar grönsaker , framförallt vitkål .
vann ni ?
jag kan inte göra det nu .
hur länge har Tom varit din pojkvän ?
oroa dig inte . han kan inte tyska .
slösa inte bort din tid .
han är förstapristagaren .
jag hade ingen aning .
köp en tandkrämstub åt mig när du är i affären .
det här tåget går mellan Tokyo och Hakata .
Tom har inget hem .
jag tycker om den här koppen .
jag skulle vilja hjälpa dig .
går han tidigt till skolan ?
du luktar illa .
det finns spårvagnar i Berlin .
jag är på sidan tre .
det finns några undantag .
när får jag komma härifrån ?
Tom bestämde sig för att ringa polisen .
jag önskar att du ringde Tom .
Tom är en gammal vän .
jag hinner inte det i morgon .
den var inte på ovanvåningen .
han vill fortfarande komma .
hur kan jag få dig att ändra dig ?
jag älskar den berättelsen .
jag skulle vilja prata med er igen .
han har en utländsk bil .
du ska alltid göra det rätta .
Tom blev utexaminerad från Harvard .
du kom tillbaka .
han är dj .
skadades någon ?
jag dricker mig aldrig full .
får jag äta den här kakan ?
han gjorde allt fotarbete .
jag trodde att Tom skulle säga hej .
här är ert kvitto .
du måste ha tålamod .
finns det en bensinmack i närheten ?
det börjar bli dags att gå hem .
han agerade snabbt och släckte elden .
du luktar gott .
tala aldrig med främlingar .
kan du inte skriva med kulspetspenna ?
har Tom barn ?
Tom är knappt vid liv .
Tom tenderar att prata ganska snabbt .
ge mig ditt sidovapen .
jag är förskräckt .
ser du den ?
jag kände mig väldigt lättad när jag hörde nyheterna .
hade du kul på turnén ?
hur klarade de sig ?
jag är trött på tv .
vad har ni hittat ?
har du något att tillägga ?
Tom och Mary vill ha vår hjälp .
Tom är eländig .
har du beställt ?
han försökte ta på sig sina nya skor .
jag måste avskeda Tom .
varför behöver du mig ?
han förstår Er inte .
han sa åt eleverna att vara tysta .
var ligger den kanadensiska ambassaden ?
de lät mig vänta länge .
jag har förfärliga nyheter .
din son är en ängel .
de är alla lika .
jag har känt henne i över 20 år .
ta en smutt av det här .
kan du ursäkta mig ?
välkommen hem till oss .
hur vet du om någon är en löpare ?
allt är annorlunda .
jag känner mig konstig idag .
också jag tycker om godis .
släpp ut mig härifrån .
de var ansvariga för olyckan .
kom prick klockan tio .
Tom tog tag i Marys hand .
jag försöker helt enkelt att inte tänka på det .
Tom blev förlägen .
jag är upprörd .
vi är föräldrar .
ni måste låta mig hjälpa till .
jag sover inte så mycket .
jag kan knappt se dig .
jag vill dricka .
Tom kände sig väldigt ensam .
vill du spela tennis med oss ?
vilket parti tillhör du ?
ge Tom lite tid .
klubben har trettio medlemmar .
varje del av ön har blivit utforskad .
hur är det relevant ?
min bror kan komma att behöva en operation för knäskadan .
varför vill du ha den här ?
byggnaden totalförstördes i jordskalvet .
han säger att hans son kan räkna till hundra nu .
jag gav dem en present på deras årsdag .
Tom är inte svag .
jag måste vara där .
lägenheten jag bor i är inte särskilt stor .
Blås ut ljusen och önska dig någonting !
våren är min favoritårstid .
jag vill träna .
det fanns ingenstans att köpa mat .
han heter Tom , inte John .
jag vill ha cashewnötter , inte mandlar .
det ligger en bok om dans på skrivbordet .
jag var tvungen att lita på Tom .
han vet bättre än att gifta sig med henne .
hur mycket kostar det där ?
kan du skilja på vete och korn ?
jag behöver en vecka .
stanna kvar .
Tom vill verkligen åka till Boston .
du verkar lycklig .
jag är inte lycklig .
jag kan inte böja min högerarm .
köpte du dem ?
är jag för krävande ?
lyssna noga !
det var söndag i går , inte lördag .
tio år har gått sedan jag kom hit .
det var väldigt roligt .
det är väldigt snällt av dig att säga det .
ingen annan än du kan göra mig lycklig .
ön ligger på ungefär två mils avstånd från kusten .
du måste vänta på nästa buss .
Tom är vänlig och givmild .
huset står i brand .
rock tilltalar unga män och kvinnor .
du måste ta tolvan .
Tom äter frukost .
jag lånade honom lite pengar , men har inte återbetalat dem än .
de krävde stränga straff för de södra rebellerna .
kan vi prata på insidan ?
var inte så negativ .
jag skulle vilja spela tennis .
han springer .
kan vi gå ut och prata ?
Räck upp handen om du vet svaret .
jag stannar här .
vad är din plan ?
när behöver Tom det ?
jag kommer känna mig ensam när du har gått .
jag visste att ni skulle vara upptagna .
sluta gnäll !
du är bedårande .
får vi vara med ?
jag kommer att vara hos Tom .
jag är glad att Tom är borta .
hur mår du ?
jag tror inte att Tom gjorde något med den .
släpp min hand .
tycker du att Tom är orättvis ?
du borde kanske skaffa en hund .
ni skrämmer mig inte .
jag gör det för att jag måste .
Tom är modfälld .
jag vill ha den där katten .
var snäll med din mamma .
jag vill åka till ett annat land .
jag gav Tom ett val .
gå före du , Tom .
kan jag ställa ned den här ?
jag förstår dig till en viss grad .
Invånarna i den här byn lever i harmoni med naturen .
du har aldrig varit bra på att rita .
choklad görs på kakaobönor .
jag avskydde det först .
vi behöver hjälp här uppe .
jag förmodade att jag skulle vara säker här .
vad har vi ?
din idiot !
jag måste hålla mig lugn .
kan du säga namnet på en av deras låtar ?
jag tar ett bad varannan dag .
var ligger närmaste museum ?
ta fram din plånbok .
ge mig min öl .
en dag kommer du att glömma bort mig .
jag går hem .
tycker du om Earl Grey @-@ te ?
otroligt , eller hur ?
minns ni den här leken ?
jag hinner inte med det i morgon .
stör det dig om jag sätter på tv:n ?
svara på frågan .
jag gick aldrig och la mig .
Tom kom fram bakom gardinen .
vi hör inget .
vår nya skolbyggnad håller på att byggas .
vill ni inte höra min version ?
Tom gjorde klart läxan innan kvällsmaten .
Tom säger att han är hungrig .
när ska du åka till Europa ?
hans tal fångade vår uppmärksamhet .
de ser honom som en hjälte .
han studerade hur fåglar flyger .
gå inte nära hunden .
var är kaptenen för det här skeppet ?
jag kan inte se något med mitt högra öga .
de två nationerna har starka affärsförbindelser .
det finns en hake .
jag tänker kasta ut Tom .
en röd klänning ser bra ut på henne .
jag älskar fjärilar .
att flyga drake kan vara farligt .
är vi klara nu ?
jag trodde att Tom var död .
jag hade en katt .
Tom tog inte självmord .
jag trodde att du var upptagen .
jag mår bra nu .
han går alltid med ett gevär i handen .
Tom Jackson blev 93 år gammal .
jag behöver den senast i morgon .
vi spelade baseball .
hur bröt du den ?
jag älskar linssoppa .
det har slutat regna .
ge mig ett val .
jag måste hem .
min fru är läkare .
jag känner mig illamående .
Tom säger att ni är bra på tennis .
ni kan inte lämna mig .
vilket språk talas i Egypten ?
jag kommer .
det går bra för Tom i skolan .
han slutade dricka .
så dyrt var det inte .
varför sa du nej ?
alltid när jag ser dig , säger mitt hjärta att jag är förälskad .
sådant händer .
spelar det någon roll ?
hur går det för mig ?
jag är studerande .
jag tror inte att kärlek finns .
han la boken på hyllan .
min bror är väldigt lång .
jag var med någon .
se till att Tom ringer mig .
du måste stanna .
vad var det i kuvertet ?
jag kunde ta en öl .
ring polisen .
min far är så att säga en vandrande ordbok .
hur gillar du stan ?
vad är klockan ?
hur mycket kostar apelsinerna ?
vad ska du göra på Halloween ?
sade Tom verkligen det ?
Tom blev fast .
Tom är fast besluten .
16 kilometer är inte en kort sträcka .
jag vet inte vad han har råkat ut för .
hon förlängde sin vistelse med fem dagar .
det kändes som om mitt ansikte brann .
det är inte något misstag .
var snäll och avbryt mig inte .
du frågar fel person .
Tom är kortare än jag .
jag sätter in tiotusen yen varje månad .
hon log åt sig själv i spegeln .
jag skulle göra vad som helst för er .
är ni tokiga ?
han är min bror .
han säger alltid ett ord för mycket .
är du rädd nu ?
Tom är driftig .
välkommen till mitt liv .
var gör det ont ?
den där simbassängen ser verkligen inbjudande ut .
minns du den här leken ?
Tom jobbar med din bil .
här kommer de .
jag avskyr karaoke .
jag ger dig mitt ord .
Tom är bara rädd .
det här var en dålig idé .
han har gått ur tiden .
de är kanske upptagna .
jag kan inte hjälpa er .
gick du i skolan i dag ?
vi kan tala med Tom .
få bort Tom härifrån .
Tom vinner .
biljetterna är slutsålda .
jag måste kolla .
vad för slags hund är det här ?
får jag äta den här tårtan ?
hans frånvaro i går berodde på förkylning .
jag gick med på att köpa den .
jag tappade tålamodet .
kan du hjälpa mig att hitta min hund ?
vi hade en underbar semester i Sverige .
Tom andas knappt .
den är noggrann .
jag håller på att bli bättre .
nu gör vi det på mitt sätt .
den här bussen får plats med femtio personer .
kan jag få mina nycklar ?
stranden är ett idealiskt ställe för att barn att leka .
Tom bestämde sig för att säga upp sig .
har Tom den ?
han tyckte inte att det var roligt .
är du min läkare ?
kaffe vore trevligt .
jag är Toms vän .
vad kommer du göra om det händer ?
Tom är Marys granne .
Fåglarna sjunger .
jag är från Ryssland .
var är Toms klassrum ?
jag har ett komplicerat ärende jag vill diskutera med dig .
ni ville att det skulle bli så här , eller hur ?
jag följde Tom dit .
eftersom så många människor vill ha ett europeiskt pass håller andelen skenäktenskap på att öka .
det här är en katastrof .
säg : &quot; kan jag få &quot; .
hämta din jacka , Tom .
jag har ingenstans att gå .
vad ska vi säga till Tom ?
han hatar spindlar .
kan du snälla säga hur lång du är och din vikt ?
Tom sade att han hoppades att du skulle vilja göra det
jag klättrade upp i ett träd .
jag vill be dig om en tjänst .
det var bara en liten kärleksaffär .
det är förmodligen hemsökt .
de såg efter pojken .
hämta mina tabletter .
vad studerade du ?
hon övertalade honom att göra det fastän hon visste att det inte var en god idé .
det är läggdags .
jag hör skratt .
pengar växer inte på träd .
kan Tom göra det ?
jag är så mätt .
Tom var tokförälskad i Mary .
jag var på bio .
hur arg är du då ?
hör du det ?
Vilka pratade ni med ?
se på alla dessa askar .
alla deltog i halloweenfesten .
jag skulle just gå .
Tom blev stor .
det doftar av blommor .
hur är det med din syster ?
förr eller senare kommer jag att slå dig .
hennes klänning var billig .
jag gick hemifrån vid sju .
jag har nyss fyllt trettio .
jag tror hur som helst inte på det .
min nätförbindelse är långsam .
stick härifrån , ungjävlar !
han har studerat utomlands .
den är god .
gå tillbaka in dit .
det är min cd @-@ skiva .
jag skjuter dig .
spara den till senare .
har du duschat ?
han gillar verkligen musik mycket .
kom och hämta mig .
kom ombord .
jag klarar inte av sådana här filmer .
Tom är handikappad .
Tom berättade för oss att det var ett gammalt skepp .
Streta inte emot .
jag sprang till min mamma .
jag lämnade Tom i sticket .
Tom visste vad han gjorde .
det finns många gamla tempel i Kyoto .
han misstar mig alltid för min syster .
hur mycket älskar du Tom ?
vi får den gratis .
jag har ett liv .
jag tror att vi har råd .
Tom berättade för Mary att John var gift .
är Ginza Japans livligaste gata ?
jag hade en blixtrande huvudvärk .
killar är dumma .
är det utegångsförbud ?
vi har ett val nu .
jag är inte färdig än .
låt mig hjälpa dig upp .
får jag ta tre ?
man kan inte lära gamla hundar sitta .
Tom är elak .
kan vi gå in och prata ?
ge mig några minuter .
jag såg Tom blinka .
du måste inte säga någonting om du inte har lust .
kan jag ställa ner den här ?
den sitter på ditt bord .
jag såg allt .
kom till festen .
lämna min familj ifred .
han blev en berömd skådespelare .
svara .
det finns ett hotell här .
efter att vi gått ett tag , kom vi fram till sjön .
jag har bara gjort detta en gång innan .
Tom råkade ta sönder sin favoritkopp .
Tom är på väg .
det är dags att stiga upp .
låt mig vara .
Tom är underhållande .
jag känner din bror ?
jag kopplade bara av .
Tom ser skamsen ut .
jag borde vila upp mig lite .
bara kärlek kan krossa ens hjärta .
du gör ett bra jobb .
män är svin .
Tom och Mary ser så lyckliga ut .
jag vill städa huset innan mina föräldrar kommer tillbaka .
vad missade vi ?
jag kommer ihåg er . vi träffades för tre år sedan .
du är inte så galen .
jag är överraskad att du vann priset .
jag tror att jag äntligen ska pensionera mig .
det är dags för tårta .
den sitter på ert skrivbord .
de hurrade .
Tom vet inte vart han skall gå .
kan ni inte se det ?
snälla gå ut härifrån genast .
det där är ett gammalt skämt .
jag ska ge dig ett exempel .
hon valde skorna som passar till klänningen .
du har spillt lite ketchup på din slips .
mördade du Tom ?
vi kan använda den .
det värsta med sommaren är hettan .
ingen kommer att beskylla dig .
jag måste få det där .
kom och träffa några av dina nya klasskamrater .
du är oansvarig .
jag behöver män som du .
Tom gillar att äta kall pizza till frukost .
vill ni inte säga någonting , behöver ni inte det .
min katt dog igår .
vi är båda mycket äldre nu .
vad har du ?
har klimatet förändrats ?
han är inte vad han utger sig för .
jag gav dig en bok .
jag är översynt .
Kortkorta kjolar har blivit omoderna .
jag måste köpa en .
har du någonsin sålt en bil ?
Tom var högt utbildad och talade åtskilliga språk flytande .
jag hoppas att det här är början på en vacker vänskap .
ge det till henne .
vi kommer att behöva ett lån .
är det någon hemma ?
jag vill ha alltihop .
jag är högerhänt .
han är irriterande .
jag tvivlar på det .
jag trodde att jag var trevlig .
jag vill lära mig standardengelska .
ta en titt på det där .
jag läste ut boken i går kväll .
är ni studenter ?
jag älskar katter också .
såg Tom dig ?
jag tog Tom till sjukhuset .
jag har ingenting att skriva med .
han blir sällan arg .
Tom lånade mig den där DVD:n .
en gång räcker inte .
hur kunde du gissa ?
jag är inte säker på när han kommer att komma .
ni verkar förvånade .
hur länge har vi på oss ?
känner du lukten av rök ?
varför är du arg på honom ?
det kommer att ordna sig .
du verkade inte förstå vad Tom sa .
byggnaden rasade samman i jordbävningen .
jag fick nästan en hjärtattack .
varför gjorde de det ?
frågade du Tom ?
målade du den här ?
jag hade en dålig natt .
han är min bror .
sa Tom när han skulle komma fram ?
hur ser du om någon är en löpare ?
