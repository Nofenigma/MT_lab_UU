kan vi gå in ?
jag är en oskyldig man .
Ryck upp dig .
Tom säger att han inte har några fiender .
Tom måste få hjälp .
ur vägen för mig .
Tom har ännu inte svarat .
ni får inte komma för sent den här gången .
jag började jobba igen .
det känns riktigt bra .
Tom är rädd för läkare .
jag är inte hungrig längre .
vi var stolta över Tom .
ät lunch med mig .
Tom är inte svag .
varför bestämde du dig för att prata om det nu ?
det där är boken som jag vill läsa .
jag läste en bok medan jag åt .
vi kommer inte att rösta på Tom .
jag är trött .
har du ätit lunch än ?
sa jag inte just det ?
jag skulle vilja tala en stund med Tom mellan fyra ögon .
han ser trött ut .
jag är ledsen , den här är inte till salu .
Tom gillar inte öl .
en sjukdom förhindrade honom från att gå ut .
Italien är inte Grekland .
gör det fort .
Tom anlände trettio minuter sen .
jag vill bara inte att Tom lägger sig i .
ge den en sekund .
gå och hämta lite verktyg .
har du fler än en mobiltelefon ?
jag måste sparka Tom .
jag skrattade mycket .
ingen kommer att klandra er .
kanske stannar jag .
Tom är tjock .
vad läser du ?
många träd tappar sina löv på vintern .
vi väntade .
hur kan du stå ut med den där killen ?
kan jag få prata med dig ?
det är inget att vara ledsen över .
ditt namn är nu borttaget från listan .
vi spelar ofta schack .
du måste få tillräckligt med sömn .
jag åt kaviar .
jag skulle vilja prata med dig igen .
många européer besöker Egypten varje år .
Olyckligtvis pratade Tom bredvid mun .
varför gör du så mot mig ?
jag är faktiskt väldigt upptagen .
han bröt reglerna .
jag måste ta ett paraply med mig .
jag var på banken .
allting måste ta slut .
vad gav Tom dig i födelsedagspresent ?
så fort det blir mörkt börjar fyrverkeriet .
varför berättade du inte det här för polisen ?
är du lärare eller student ?
Tom alltid på sig en hatt .
kan vi inte bara spankulera runt i parken ?
jag kan hämta den .
Tom har bestämt sig för att klippa sig först till våren .
Toms katt fick nio kattungar .
jag borde aldrig ha sagt mitt lösenord till Tom .
Tom tog av sig skjortan .
vad finns i den här lådan ?
hur gör Tom det här ?
vad är syftet med den ?
Krokodiler har vassa tänder .
jag glömde min jacka .
det stämmer !
han är österrikare .
Tom är en hippie .
jag var inte skyldig Tom någonting .
du är tillräckligt gammal för att förstå .
har den ett badrum ?
jag tycker verkligen om det .
hans föräldrar älskar mig .
Tom räddade mig .
jag är mjuk i lederna som en akrobat .
Tom sköljde schampot ur sitt hår .
jag tänker inte diska .
vem hatar er ?
Tom högg Mary i nacken med sin kulspetspenna .
jag har väldigt ont .
jag är elev .
det är molnigt .
Tom är motbjudande .
skolan ligger en halv mils promenad från mitt hus .
Tom försvann snabbt i vimlet .
han är lika lång som min far .
god morgon .
vet du vilken färg hon tycker om ?
jag vill ha ett eget rum .
vi åt lunch .
det kan komma att göra ont .
håll ut , Tom .
Tom gick precis in .
vänta tills sex .
Tom hatar insekter .
jag hatade det i början .
ni är farliga .
jag ska försöka att fixa det här , men det kan hända att jag inte lyckas .
han stoppade näsduken i sin ficka .
när jag hittade rummet var det tomt .
Kanada producerar bra vete .
Tom sparkade omkull en stol .
vi associerar Egypten med Nilen .
jag tycker att Tom är ambitiös .
har Tom fått sparken än ?
jag har rätt att vara på det här skeppet .
ta god tid på dig .
Grytan var min .
jag vet inte när jag kommer att kunna hjälpa dig .
lova mig att inte skratta .
jag arbetar 3 timmar varje söndagsmorgon .
jag trodde att fienden hade dödat Tom .
Solenergi är miljövänlig .
jag är här för att anmäla ett brott .
hur gick det på jobbet ?
hur länge sen är det ?
har du designat den här ?
vad gjorde Tom här ?
var är min tidning ?
jag kan ta hand om Tom .
klockan är 9.15 .
jag ville bara att du skulle titta på detta .
vi tog en taxi .
titta på hajarna .
jag har andra planer .
min kropp är inte så smidig som den brukade vara .
en dag kommer ni att ångra det här .
du är en bra tennisspelare .
Ställ er upp , allesamman .
det var fullmåne i går .
det betydde mycket för mig .
jag har nariga läppar .
jag vill drömma .
jag tycker att du borde berätta för Tom att du älskar honom .
jag är lycklig här .
Tom sade åt Mary att ljuga .
jag tänker så det knakar , men jag kan inte komma på hennes namn .
Tom är tveksam .
du borde stanna .
jag är glad att vi gjorde det där .
de ser alla lyckliga ut .
det är en slags katt .
hur länge kommer det här kalla vädret att hålla på ?
han gick och lade sig klockan tio som vanligt .
förlät Tom dig ?
jag är glad att Tom ska hjälpa oss .
måste jag betala dig ?
förresten , spelar du fiol ?
jag gick inte , utan stannade hemma .
kan ni reparera detta ?
ursäkta mig en sekund .
det är någonting som inte stämmer här .
ett enormt monster är på väg ned från berget .
jag spelar gitarr .
jag är inte intresserad .
jag såg matchen .
du har två kulor .
får jag träffa Tom idag ?
jag är er advokat .
var lärde ni er att skriva ?
använd den här .
vi välkomnar alla som vill komma till festen .
är era väskor packade ?
jag ångrar det inte alls .
jag har aldrig hört talas om er .
Dinosaurierna dog ut för en mycket lång tid sedan .
detta är riktigt illa .
jag lade märke till att hon satt på främsta raden .
jag kommer inte att vänta för alltid .
jag köpte en sax .
det är en risk som Tom måste ta .
jag ska spela fotboll efter skolan .
ursäkta , kan du förklara vägen till stationen ?
det är min hemlighet .
jag ska till Paris i helgen .
Tom och Mary paddlade kanot längs med floden sist jag såg dem .
ge den ett ögonblick .
jag har inte på mig den här .
Tom är ursinnig .
Tom hatar oliver .
stäng igen er bok .
ta reda på var Tom är .
det kan inte vara så dåligt .
jag är vid den norra utgången .
jag gav Tom trettio dollar .
vi kommer att behöva Toms hjälp .
ikväll ska jag stanna hemma .
det är ingen hemlighet .
följde någon efter oss hit ?
jag känner till det .
jag klippte mig i fingret .
var hänsynslösa .
jag träffade Tom några veckor innan han dog .
jobbar de här ?
det är bäst att du inte väntar längre .
så romantiskt !
jag tappade bort min anteckningsbok .
den är inte klar än .
hon kysste honom på pannan .
jag var vacker en gång .
regnet slog emot fönstren .
ni måste inte komma hit varje dag .
träffade du Tom ?
min fråga är varför .
jag håller på att bli galen .
är det inte bättre så här ?
vill du ha lite öl ?
Åk till sjukhuset .
de var falska .
en minderårig är beroende av sina föräldrar .
Tom saknas .
jag är i bilen .
jag matade hunden .
jag skulle vilja äta frukost med dig .
vi turades om att köra .
jag klandrar dig inte det minsta .
någonting är inte rätt här .
tittar de på oss ?
det snöar i Paris .
om du vill ha fred , förbered dig för krig .
de jobbar på övervåningen .
jag utmanar dig på tennis .
hur kan vi hjälpa till ?
vad köpte Tom till dig ?
kan någon bevisa det ?
när såg du henne senast ?
jag ska ta min rock .
de kommer att ha jättekul .
jag träffade ingen på vägen hem .
jag trodde att det var ett skämt .
jag tror att Tom hade rätt .
behöver jag någon medicin ?
hur säger du det på italienska ?
jag önskar att jag hade en bil .
jag stavade ordet fel .
kan vi lita på dem ?
blev du rånad ?
jag ger mig av nu .
kom tillbaka !
jag är säker att Tom inte kommer hålla med
det är precis vad Tom behöver .
jag var närvarande i skolan igår .
alla pojkarna sprang iväg .
jag kan inte bekräfta det .
jag trodde att du gick hem .
var vänlig , men bestämd .
jag tycker bättre om dig .
jag köpte den här åt dig .
jag är nöjd här .
jag har goda nyheter .
tycker du om ost ?
Tom är skild .
hur mycket kostade det ?
han har alltid för lite pengar .
vanligtvis kan Tom få vad han vill .
Tom gav ett ben till sin hund .
ät så mycket du vill .
Tom visste att jag var redo .
jag fick ge upp .
jag kan föra dig dit .
jag antar att det inte är så enkelt .
hur kan vi hjälpa till ?
jag kan inte göra det här .
jag tänker inte hindra dig .
han är bara en vanlig kontorsråtta .
jag gav inte Tom något val .
du är singel , eller hur ?
på vems sida är ni ?
jag gjorde det inte .
det här är den högsta byggnad som jag någonsin har sett .
jag kommer tillbaka om 2 veckor .
var det inte rödvin du beställde ?
vi kommer inte att kunna ringa dig .
hon kysste honom .
vet ni ens vem Tom är ?
Tom kan ännu vara vid liv .
jag har jobbat med det här i tre veckor .
hur återhämtar man sig från någonting sådant ?
katten är på mattan .
man ska inte döma folk efter utseendet .
vi förlorade .
är du redo för att lära dig sanningen ?
spelet är inte över .
många människor litar inte på regeringen .
vad innebar det ?
kan du gå , Tom ?
jag vet hur mycket du älskar Tom .
jag är tacksam för er hjälp .
vi gick redan igenom det där .
jag har inte bestämt mig än .
släpp min son .
jag hittar inte min portfölj .
när börjar vi ?
känner ni dem ?
det var en stor en .
Tom är en väldigt dålig kille .
hans fru är en synnerligen begåvad kvinna .
hur lång tid har du på dig ?
Tom är fortfarande vaken .
det här är skandalöst !
jag lagar mat .
den här skulpturen är mer än två tusen år gammal .
vad vill du då ?
jag har gömt den någonstans .
allt är normalt .
han har redan gått .
jag var artig .
jag skulle vilja följa med Tom .
jag kan vänta .
jag vill färga mitt hår rött .
det har varit mulet de senaste dagarna .
är du nästan framme ?
du bör följa skolans regler .
lämna mig i fred .
var snäll och säg svaret på frågan .
jag hoppas att jag vinner .
är det där Tom ?
han studerar alltid flitigt .
jag planerar att ge min son en dator i slutet av månaden .
Tom bodde på övre våningen .
det är apkött .
stal du den här ?
snabba er , ungar , annars missar ni skolbussen .
jag har en båt och en bil .
ingenting spelar egentligen någon roll .
har du sovit ?
planet har nyss lyft .
jag ska göra det för dig .
Tom gjorde mål .
jag kan inte göra detta utan er .
vad smart !
det är något med honom som jag inte gillar .
de avisade bron med salt .
de flesta amerikanare tycker om hamburgare .
jag litar på dig .
ring mig senare .
jag älskade verkligen Tom .
jag önskar att jag ringt Tom .
jag tycker om att spela tennis och golf .
ser ni någonting ?
&quot; han har varit sjuk &quot; . &quot; Jaså , jag hoppas att det inte är någonting allvarligt &quot; .
Tom är den enda jag känner som kan göra det här .
de simmade ut till ön .
jag vill inte spela .
jag tycker det här vinet är bra .
var ska vi ses ?
snälla , lämna oss inte här .
det kommer inte att göra ont .
kolla det här .
ni kunde ha dött .
Tom är sjuk .
jag sa det till Tom själv .
jag vet vad som är fel .
hur många tog du ?
jag håller ett säte åt dig .
jag måste fokusera .
det röda paraplyet påminde henne om hennes farmor .
han är en man som man kan räkna med .
Tom ser sjuk ut .
Tom höll med om allting Mary sa .
vi ska göra det igen .
sätt er .
jag blöder om knät .
Tom är en tävlingsmänniska .
jag vill bara vila .
vad är er fars namn ?
Tom är vanvettig .
jag förstår mig inte på honom .
ha en trevlig flygresa .
det röda paraplyet påminde henne om hennes mormor .
Vilka vill ni tala med ?
Körsbär är röda .
jag gjorde dig en tjänst .
vi har diskuterat det här problemet nyligen .
jag vill sova .
Tom kallade Mary för dumbom .
vad har jag missat ?
bli inte stött . Tom är så där med alla .
ta en karta med dig ifall du skulle gå vilse .
Hotar du mig ?
Fortsätt söka .
ni borde vara försiktigare nästa gång .
gå inte ut på framsidan .
hämta min mat .
hon gillade poesi och musik .
alla tittade .
jag är en lycklig man .
hans chef är väldigt krävande .
kan jag få ett glas vatten , tack .
det där är min pappa .
vi vill bara ha dig .
sylt fås på burk .
jag gillar den där klänningen .
har du fördomar ?
kan du göra det eller inte ?
vilken är din favoritsaga ?
jag har varit med om en olyckshändelse .
jag såg slagsmålet .
jag är bara en taxichaufför .
gör som ni vill .
jag glömde att låsa ytterdörren .
vi måste vänta och se .
det här kan vara ett undantag .
Välj ett lösenord som är lätt att komma ihåg , men svårt att gissa sig till .
jag bor inte i Boston .
hur många hästar äger Tom ?
Tom kunde inte bryta sig in i den .
jag sa åt Tom att han inte skulle komma idag .
här är hon !
ta det lugnt .
dagarna blir längre och längre .
följer du efter mig ?
hur mår din pappa ?
jag vet att ni saknar er familj .
jag tycker om att mata duvorna .
köpte du Tom en hund ?
jag var förälskad .
jag kan ringa Tom .
jag röstade inte på någon .
Tom visste inte vad Mary planerade .
jag förtjänar inte att leva .
vilken är nästa station ?
det är inte så litet .
hur tog du dig hit ?
tala i mikrofonen .
Basketlaget tränar inte på måndagar .
han bakade muffins .
det var ingen jordbävning .
vad har du för order ?
ingen sprang före honom .
vad viskar du för ?
Sväng vänster .
det landet har ett handelsöverskott . det exporterar mera än det importerar .
Tom visste att jag var på väg .
när startar vi ?
reglerna är inte viktiga .
jag ska ta hand om det .
jag var där först .
ni har vuxit .
jag ville inte skryta .
är du fortfarande hungrig ?
jag bryr mig inte om vad Tom gör .
de ringde .
jag lyssnar på musik .
hon hittade jobb som maskinskriverska .
de har ingen annanstans att gå .
ett äpple om dagen håller doktorn borta .
det måste finnas ett mönster .
var allvarlig .
jag tycker om godis också .
tänker du på franska ?
hade jag något val ?
han har ingen dator .
Tom sa att han ville dö .
sluta göra omsvep och kom till saken .
Tom gav Mary en kopp .
jag tycker bättre om grapefrukter än apelsiner .
jag är lite tokig .
jag skulle vilja stanna så länge som möjligt .
Tom såg videon .
varför hatar du Tom ?
Tom blev tvungen att improvisera .
det sker automatiskt .
mitt flyg var inställt .
den måste tas bort .
jag vill egentligen bara skaffa vänner .
ringde Tom ?
kan ni höra mig ?
vill du ha en banan ?
Fåglarna flög söderut .
jag är lite hungrig .
jag är ingen profet .
Tom har erkänt .
det finns ingenting du kan göra .
kan du säga det en gång till ?
de kör fast .
du verkar vara förvånad .
Tom skäms .
jag vill ha det där jobbet .
hur går det med skolan ?
han vill inte vänta på dig .
hur mycket vill du ha ?
allt är okej .
vad kostar det här paraplyet ?
min far insisterade på att vi skulle vänta på tåget .
vad var problemet ?
vad kan du se ?
är den vit ?
jag vill ha mera mjölk .
hur överlevde Tom ?
jag ska gå och fråga Tom .
